(0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")),
1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14|15|16|21|22|23|24 => Pixel_t'("00","01","00"), 17|18|19|20 => Pixel_t'("01","01","01")),
2 => (0|1|2|3|4|5|6|7|8|9|10|11|12|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 13|23 => Pixel_t'("00","01","00"), 15|16 => Pixel_t'("00","01","01"), 14 => Pixel_t'("01","01","01"), 21|22 => Pixel_t'("01","10","01"), 17|20 => Pixel_t'("01","10","10"), 18|19 => Pixel_t'("10","11","10")),
3 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17 => Pixel_t'("01","01","01"), 22|24 => Pixel_t'("01","10","01"), 21 => Pixel_t'("01","10","10"), 19|20|23 => Pixel_t'("01","11","10"), 18 => Pixel_t'("10","11","10")),
4 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 23|25 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 18|19|24 => Pixel_t'("10","11","10")),
5 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","10","01"), 26 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 19|23|24|25 => Pixel_t'("10","11","10")),
6 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 28 => Pixel_t'("00","01","00"), 25 => Pixel_t'("01","10","01"), 26|27 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 19|23|24 => Pixel_t'("10","11","10")),
7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","01","00"), 26 => Pixel_t'("01","10","01"), 27 => Pixel_t'("01","10","10"), 21|24|25|28 => Pixel_t'("01","11","10"), 19 => Pixel_t'("10","10","10"), 20|22|23 => Pixel_t'("10","11","10")),
8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 30 => Pixel_t'("00","01","00"), 19|25|26|27|28|29 => Pixel_t'("01","10","01"), 21|22|23|24 => Pixel_t'("01","11","10"), 20 => Pixel_t'("10","11","10")),
9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 31 => Pixel_t'("00","01","00"), 19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'("01","10","01")),
10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 22|26|32 => Pixel_t'("00","01","00"), 21 => Pixel_t'("00","01","01"), 19|23|24|25|27|28|29 => Pixel_t'("00","10","01"), 17|18|20|30|31 => Pixel_t'("01","10","01")),
11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 16|19|20|21|23|26|27 => Pixel_t'("00","01","00"), 22|24|25 => Pixel_t'("00","10","00"), 28|29|30|31 => Pixel_t'("00","10","01"), 17|18|32 => Pixel_t'("01","10","01")),
12 => (0|1|2|3|4|5|6|8|9|10|11|12|13|14|15|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 7|16|18|19|20|21|23|24|25|27|28|29|32|33 => Pixel_t'("00","01","00"), 31 => Pixel_t'("00","01","01"), 22 => Pixel_t'("00","10","00"), 26|30 => Pixel_t'("00","10","01"), 17 => Pixel_t'("01","10","01")),
13 => (0|1|2|11|12|13|14|15|36|37|38|39 => Pixel_t'("00","00","00"), 3|4|9|10|16|28|29|32 => Pixel_t'("00","01","00"), 35 => Pixel_t'("00","01","01"), 27 => Pixel_t'("00","10","00"), 5|6|7|8|18|19|20|25|26|30|31|33 => Pixel_t'("00","10","01"), 17|21|22|23|24|34 => Pixel_t'("01","10","01")),
14 => (0|1|9|10|39 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|11|13|29|30|31|32|33|34|35|36|37|38 => Pixel_t'("00","01","00"), 12 => Pixel_t'("00","01","01"), 14|15|26|27|28 => Pixel_t'("00","10","01"), 16|17|22|25 => Pixel_t'("01","10","01"), 21 => Pixel_t'("01","10","10"), 18|19|23|24 => Pixel_t'("01","11","10"), 20 => Pixel_t'("10","10","10")),
15 => (0|1|3|10|11|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 2|4|5|6|7|8|9|12|13|14|15|23|24|25|26|27|28|29|30|31|35 => Pixel_t'("00","01","00"), 16|21 => Pixel_t'("00","10","01"), 17|18|19|20|22 => Pixel_t'("01","10","01")),
16 => (0|1|2|3|9|10|11|12|13|14|15|16|32|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|5|6|7|8|21|22|23|24|25|26|27|28|29|30|31|33|34 => Pixel_t'("00","01","00"), 20 => Pixel_t'("00","10","00"), 19 => Pixel_t'("00","10","01"), 17|18 => Pixel_t'("01","10","01")),
17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'("00","01","00"), 17|18|19 => Pixel_t'("00","10","01")),
18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 16|20|21|22|23|24|25|26|27|28|29|30|31|32 => Pixel_t'("00","01","00"), 19 => Pixel_t'("00","10","00"), 18 => Pixel_t'("01","10","01"), 17 => Pixel_t'("01","11","01")),
19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28|29|30|31 => Pixel_t'("00","01","00"), 17|18 => Pixel_t'("01","10","01")),
20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18|19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'("00","01","00")),
21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","01","00")),
22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28 => Pixel_t'("00","01","00")),
23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27 => Pixel_t'("00","01","00")),
24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25 => Pixel_t'("00","01","00"), 26 => Pixel_t'("00","10","01")),
25 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25 => Pixel_t'("00","01","00")),
26 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18|19|21|22|23|24 => Pixel_t'("00","01","00"), 20 => Pixel_t'("00","10","01")),
27 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17|18|19|22|23 => Pixel_t'("00","01","00"), 14|21 => Pixel_t'("00","01","01"), 20 => Pixel_t'("00","10","01"), 15|16 => Pixel_t'("01","01","01")),
28 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|22|23|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17|24 => Pixel_t'("00","01","00"), 14|15|16|18|21 => Pixel_t'("00","01","01"), 19|20 => Pixel_t'("01","01","01")),
29 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")));