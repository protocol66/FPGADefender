(0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00")),
1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|26|27|28|29 => Pixel_t'("00","00","00"), 16|23|24 => Pixel_t'("00","01","00"), 19 => Pixel_t'("00","01","01"), 18|20|21|22|25 => Pixel_t'("01","01","01"), 17 => Pixel_t'("01","10","10")),
2 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("00","01","00"), 14 => Pixel_t'("01","01","00"), 16|17|18|19|20|21|22|23|24 => Pixel_t'("01","01","01"), 25 => Pixel_t'("10","10","10")),
3 => (0|1|2|3|4|5|6|7|8|9|10|11|12|27|28|29 => Pixel_t'("00","00","00"), 13|15|16|17 => Pixel_t'("00","01","00"), 24 => Pixel_t'("00","01","01"), 18|19|20|21|22|23|26 => Pixel_t'("01","01","01"), 14 => Pixel_t'("01","10","01"), 25 => Pixel_t'("10","10","10")),
4 => (0|1|2|7|8|9|10|11|12|18|19|20|21|22|29 => Pixel_t'("00","00","00"), 3|4|6|16|17|23|24 => Pixel_t'("00","01","00"), 5|13|26|27|28 => Pixel_t'("01","01","01"), 14|15 => Pixel_t'("01","10","01"), 25 => Pixel_t'("01","10","10")),
5 => (0|1|18|19|20|21|22 => Pixel_t'("00","00","00"), 9|12|13|14|15|16|17|23|24|26|27 => Pixel_t'("00","01","00"), 2|3 => Pixel_t'("01","01","00"), 4|8|10|11|29 => Pixel_t'("01","01","01"), 5|6|7|25|28 => Pixel_t'("01","10","01")),
6 => (0|14|15|19|20|21|22 => Pixel_t'("00","00","00"), 1|2|3|12|13|16|17|18|29 => Pixel_t'("00","01","00"), 4|5 => Pixel_t'("01","01","00"), 6|7|8|9|11|23|24|25|26|27|28 => Pixel_t'("01","01","01"), 10 => Pixel_t'("01","10","01")),
7 => (0|1|29 => Pixel_t'("00","00","00"), 2|3|4|5|7|8|9|10|11|12|13|14|15|16|17|28 => Pixel_t'("00","01","00"), 18|19 => Pixel_t'("01","01","01"), 6|20|22|25|26|27 => Pixel_t'("01","10","01"), 21|24 => Pixel_t'("01","10","10"), 23 => Pixel_t'("10","10","10")),
8 => (0|1|2|3|4|5|7|8|9|10|11|12|13|14|15|16|28|29 => Pixel_t'("00","00","00"), 6|17 => Pixel_t'("00","01","00"), 27 => Pixel_t'("01","01","01"), 18|19|26 => Pixel_t'("01","10","01"), 20|21|23 => Pixel_t'("01","10","10"), 22|24|25 => Pixel_t'("10","10","10")),
9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|27|28|29 => Pixel_t'("00","00","00"), 26 => Pixel_t'("01","01","01"), 17|18 => Pixel_t'("01","10","01"), 19|20|21|25 => Pixel_t'("01","10","10"), 22|23|24 => Pixel_t'("10","10","10")),
10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|25|26|27|28|29 => Pixel_t'("00","00","00"), 16|24 => Pixel_t'("01","01","01"), 17 => Pixel_t'("01","10","01"), 18|19|20|21|23 => Pixel_t'("01","10","10"), 22 => Pixel_t'("10","10","10")),
11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 22 => Pixel_t'("01","01","01"), 16|17 => Pixel_t'("01","10","01"), 18 => Pixel_t'("01","10","10"), 19|20|21 => Pixel_t'("10","10","10")),
12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("00","01","00"), 16|17 => Pixel_t'("01","01","01"), 18|20 => Pixel_t'("01","10","01"), 19 => Pixel_t'("10","10","10")),
13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15|17|18 => Pixel_t'("01","01","01"), 16 => Pixel_t'("01","10","01")),
14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","01","01"), 15|16|17 => Pixel_t'("01","10","01")),
15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14 => Pixel_t'("00","01","00"), 18 => Pixel_t'("01","01","01"), 15|16|17 => Pixel_t'("01","10","01")),
16 => (0|1|2|3|4|5|6|7|8|9|10|11|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 12 => Pixel_t'("00","01","00"), 13|17 => Pixel_t'("01","01","01"), 14|15|16 => Pixel_t'("01","10","01")),
17 => (0|1|2|3|4|5|6|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14|15|17 => Pixel_t'("00","01","00"), 7|12|13|16 => Pixel_t'("01","01","01"), 8|9|10|11 => Pixel_t'("10","10","10")),
18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14|17 => Pixel_t'("00","01","00"), 15 => Pixel_t'("01","10","01"), 16 => Pixel_t'("10","10","10")),
19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|17|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","10","10")));