../../components/counter.vhdl