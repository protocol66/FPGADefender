library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.my_data_types.all;

package bitmaps is
    constant BACKGROUND : Pixel_t := BLACK;
    constant MAIN_CLK_FREQ : integer := 50000000;

    constant screen_HEIGHT : positive := 479;
    constant screen_WIDTH : positive := 639;

    constant pepe_sizeX : positive := 100;
    constant pepe_sizeY : positive := 100;

    constant line_sizeX : positive := screen_WIDTH;
    constant line_sizeY : positive := 2;

    constant ship_sizeX : positive := 25;
    constant ship_sizeY : positive := 25;
    
    constant laser_sizeX : positive := ship_sizeX;
    constant laser_sizeY : positive := 1;

    constant score_sizeX : positive := 15;
    constant score_sizeY : positive := 25;
    constant score_space_size :positive := 5;
    constant score_board_sizeX : positive := (score_sizeX + score_space_size)*5 + score_sizeY;
    constant score_board_sizeY : positive := score_sizeY;

    constant alien1_sizeX : positive := 20;
    constant alien1_sizeY : positive := 20;

    constant H_LINE : bit_map_t (0 to line_sizeY-1, 0 to line_sizeX-1) := (others => (others => WHITE));
    constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) := (others => (others => TEAL));
    constant LASER : bit_map_t (0 to laser_sizeY-1, 0 to laser_sizeX-1) := (others => (others => GREEN));
    constant ALIEN_1 : bit_map_t (0 to alien1_sizeY-1, 0 to alien1_sizeX-1) := (others => (others => YELLOW)); 


    constant fx1 : Sound_FX_t := (18, (550, 404, 315, 494, 182, 260, 455, 387, 340, 550, 404, 315, 494, 182, 260, 455, 387, 340, others => 0));
    constant fx2 : Sound_FX_t := (10, (300, 350, 500, 700, 990, 970, 1050, 1010, 950, 800, 770, 640, 500, 350, 355, others => 0));
    constant fx3 : Sound_FX_t := (6,  (500, 790, 950, 1300, 1710, 1650, 1300, 800, 700, others=> 0));
    constant fx4 : Sound_FX_t := (60, (1300, 1650, 1660, 1510, 1309, 1158, 1007, 855, others=> 0));
    constant fx5 : Sound_FX_t := (25, (300, 210, 310, 170, 250, 210, 310, 120, 220, 170, 160, 90, 290, 230, 140, 320, 200, 100, 250, 290, others => 0));
    constant fx6 : Sound_FX_t := (15, (700, 702, 698, 701, 699, 700, 250, 251, 249, 252, 248, 130, 131, 129, 132, 128, 130, 130, others=>0));

    constant score_9 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    constant score_8 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    constant score_7 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    constant score_6 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    constant score_5 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => PURPLE));
    constant score_4 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => YELLOW));
    constant score_3 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    constant score_2 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    constant score_1 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    constant score_0 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    constant score_blank : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BACKGROUND));
    
    -- DONT USE THIS... adds 30+ min to compile time...
    -- constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) :=
    -- (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")),
    -- 1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")),
    -- 2 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 1|2|3|4 => Pixel_t'(X"1",X"1",X"1"), 5|57 => Pixel_t'(X"2",X"2",X"2"), 54 => Pixel_t'(X"3",X"3",X"3"), 55 => Pixel_t'(X"3",X"4",X"4"), 6|36 => Pixel_t'(X"5",X"5",X"6"), 56 => Pixel_t'(X"5",X"6",X"6"), 11|12|13|14|15|31|32|33|34 => Pixel_t'(X"6",X"7",X"7"), 7|8|9|10|16|35 => Pixel_t'(X"7",X"7",X"7"), 19|20|22|24|25 => Pixel_t'(X"7",X"7",X"8"), 17|18|21|23|26|27|28|29|30 => Pixel_t'(X"7",X"8",X"8")),
    -- 3 => (38|39|40|41|42|43|44|45|46|47|48|49|50|51|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 0|37|52 => Pixel_t'(X"1",X"1",X"1"), 58 => Pixel_t'(X"2",X"2",X"2"), 53 => Pixel_t'(X"3",X"3",X"3"), 21|22|23|29 => Pixel_t'(X"6",X"6",X"6"), 19|20|24|25|26|28 => Pixel_t'(X"6",X"6",X"7"), 17|18|27 => Pixel_t'(X"6",X"7",X"7"), 1|16|32 => Pixel_t'(X"7",X"7",X"7"), 15 => Pixel_t'(X"7",X"7",X"8"), 14|30|54 => Pixel_t'(X"7",X"8",X"8"), 2 => Pixel_t'(X"8",X"8",X"8"), 4|5|13|31|33|34|35 => Pixel_t'(X"8",X"8",X"9"), 3|36|55|57 => Pixel_t'(X"8",X"9",X"9"), 12 => Pixel_t'(X"9",X"9",X"a"), 6|56 => Pixel_t'(X"9",X"a",X"a"), 7|8 => Pixel_t'(X"a",X"a",X"b"), 11 => Pixel_t'(X"b",X"b",X"c"), 9 => Pixel_t'(X"b",X"c",X"c"), 10 => Pixel_t'(X"c",X"d",X"d")),
    -- 4 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 20|21|23|26|27|28 => Pixel_t'(X"1",X"1",X"1"), 16|17|18|19|22|24|25 => Pixel_t'(X"1",X"1",X"2"), 12|13|14|15|32|51 => Pixel_t'(X"2",X"2",X"2"), 1|29|59 => Pixel_t'(X"3",X"3",X"3"), 11 => Pixel_t'(X"4",X"4",X"4"), 33 => Pixel_t'(X"5",X"5",X"6"), 31|36|52 => Pixel_t'(X"5",X"6",X"6"), 5 => Pixel_t'(X"6",X"6",X"7"), 2|30 => Pixel_t'(X"6",X"7",X"7"), 55 => Pixel_t'(X"7",X"7",X"7"), 3|4|34|35|53|54|56|58 => Pixel_t'(X"7",X"8",X"8"), 6 => Pixel_t'(X"8",X"8",X"9"), 57 => Pixel_t'(X"8",X"9",X"9"), 7 => Pixel_t'(X"9",X"9",X"9"), 8 => Pixel_t'(X"9",X"a",X"a"), 10 => Pixel_t'(X"a",X"b",X"b"), 9 => Pixel_t'(X"c",X"d",X"d")),
    -- 5 => (0|1|37|38|39|40|41|42|43|44|45|46|47|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 48|63 => Pixel_t'(X"1",X"1",X"1"), 36|49|62 => Pixel_t'(X"2",X"2",X"2"), 21|22|23 => Pixel_t'(X"2",X"3",X"3"), 16|17|18|19|20|24|25|26|27|28 => Pixel_t'(X"3",X"3",X"3"), 15 => Pixel_t'(X"3",X"3",X"4"), 14 => Pixel_t'(X"3",X"4",X"4"), 2|13|32|61 => Pixel_t'(X"4",X"4",X"4"), 12|31 => Pixel_t'(X"4",X"4",X"5"), 50 => Pixel_t'(X"4",X"5",X"5"), 3|11|29 => Pixel_t'(X"5",X"6",X"6"), 30 => Pixel_t'(X"6",X"6",X"6"), 51|60 => Pixel_t'(X"6",X"7",X"7"), 4|5|33|52|55 => Pixel_t'(X"7",X"7",X"7"), 6|10|53|54 => Pixel_t'(X"7",X"7",X"8"), 7|9|34|35|56|59 => Pixel_t'(X"7",X"8",X"8"), 8 => Pixel_t'(X"8",X"8",X"8"), 58 => Pixel_t'(X"8",X"9",X"9"), 57 => Pixel_t'(X"9",X"a",X"a")),
    -- 6 => (0|1|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 2 => Pixel_t'(X"0",X"1",X"0"), 6|7|8|9|72 => Pixel_t'(X"1",X"1",X"1"), 68|69|70|71 => Pixel_t'(X"2",X"2",X"2"), 5 => Pixel_t'(X"2",X"2",X"3"), 10 => Pixel_t'(X"2",X"3",X"3"), 44|67 => Pixel_t'(X"3",X"3",X"3"), 4|45 => Pixel_t'(X"3",X"4",X"4"), 29|30|31|32|66 => Pixel_t'(X"4",X"4",X"4"), 15|16 => Pixel_t'(X"4",X"4",X"5"), 3|11|14|33|34|43|46 => Pixel_t'(X"4",X"5",X"5"), 38 => Pixel_t'(X"4",X"7",X"8"), 12|13|19|20|21|22|23|24|28|35|40 => Pixel_t'(X"5",X"5",X"5"), 25|65 => Pixel_t'(X"5",X"5",X"6"), 17|18|26|27|41|47 => Pixel_t'(X"5",X"6",X"6"), 42 => Pixel_t'(X"5",X"7",X"7"), 39 => Pixel_t'(X"6",X"6",X"6"), 48|51|52|53|54|55|56|57|58|64 => Pixel_t'(X"6",X"7",X"7"), 49|50|59|63 => Pixel_t'(X"7",X"7",X"7"), 60|61|62 => Pixel_t'(X"7",X"8",X"8")),
    -- 7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|29|30|31|32|33|34|35|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 17|28 => Pixel_t'(X"2",X"2",X"2"), 18|19|26|43 => Pixel_t'(X"3",X"3",X"3"), 44 => Pixel_t'(X"3",X"3",X"4"), 25|27|42|45 => Pixel_t'(X"3",X"4",X"4"), 38 => Pixel_t'(X"3",X"6",X"6"), 20 => Pixel_t'(X"4",X"4",X"4"), 46 => Pixel_t'(X"4",X"4",X"5"), 21|22|24|41|47|48|49 => Pixel_t'(X"4",X"5",X"5"), 23 => Pixel_t'(X"5",X"5",X"5"), 53 => Pixel_t'(X"5",X"5",X"6"), 50|51|52|54|55|57 => Pixel_t'(X"5",X"6",X"6"), 56 => Pixel_t'(X"6",X"6",X"6"), 58|72 => Pixel_t'(X"6",X"6",X"7"), 59 => Pixel_t'(X"7",X"7",X"8"), 39|40|60|61|62|68|71 => Pixel_t'(X"7",X"8",X"8"), 69|70 => Pixel_t'(X"8",X"8",X"9"), 63|64|67 => Pixel_t'(X"8",X"9",X"9"), 65|66 => Pixel_t'(X"8",X"9",X"a")),
    -- 8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|27|28|29|30|31|32|33|34|35|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 26 => Pixel_t'(X"0",X"1",X"0"), 20|38 => Pixel_t'(X"1",X"1",X"1"), 50|51|52 => Pixel_t'(X"2",X"2",X"2"), 68 => Pixel_t'(X"2",X"3",X"3"), 21|49|53|64|65|66|67|69|70|71|72 => Pixel_t'(X"3",X"3",X"3"), 63 => Pixel_t'(X"3",X"3",X"4"), 25|59|60 => Pixel_t'(X"3",X"4",X"4"), 22|23|54|57|58|61|62 => Pixel_t'(X"4",X"4",X"4"), 55 => Pixel_t'(X"4",X"5",X"4"), 24|48|56 => Pixel_t'(X"4",X"5",X"5"), 42|45|46|47 => Pixel_t'(X"5",X"6",X"6"), 43|44 => Pixel_t'(X"6",X"6",X"6"), 39 => Pixel_t'(X"6",X"7",X"6"), 40|41 => Pixel_t'(X"7",X"8",X"8")),
    -- 9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|28|29|30|31|32|33|34|35|36|50|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 49 => Pixel_t'(X"0",X"1",X"1"), 21|27|37|48|51|52|53|61 => Pixel_t'(X"1",X"1",X"1"), 22|23 => Pixel_t'(X"2",X"2",X"2"), 58|59|60 => Pixel_t'(X"3",X"3",X"3"), 24 => Pixel_t'(X"3",X"4",X"4"), 26|54 => Pixel_t'(X"4",X"4",X"4"), 25 => Pixel_t'(X"4",X"5",X"5"), 47|57 => Pixel_t'(X"5",X"5",X"5"), 38 => Pixel_t'(X"7",X"8",X"8"), 55|56 => Pixel_t'(X"8",X"8",X"8"), 39|45|46 => Pixel_t'(X"8",X"9",X"9"), 42 => Pixel_t'(X"8",X"a",X"9"), 44 => Pixel_t'(X"9",X"a",X"a"), 43 => Pixel_t'(X"a",X"a",X"a"), 40|41 => Pixel_t'(X"c",X"d",X"d")),
    -- 10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|29|30|31|32|33|34|35|36|47|48|49|50|51|52|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 24|53|59 => Pixel_t'(X"1",X"1",X"1"), 28 => Pixel_t'(X"1",X"2",X"2"), 54 => Pixel_t'(X"2",X"2",X"2"), 25 => Pixel_t'(X"3",X"4",X"4"), 46|57|58 => Pixel_t'(X"4",X"4",X"4"), 27 => Pixel_t'(X"4",X"5",X"5"), 26 => Pixel_t'(X"5",X"5",X"5"), 37|55 => Pixel_t'(X"7",X"8",X"8"), 45 => Pixel_t'(X"8",X"8",X"8"), 56 => Pixel_t'(X"8",X"9",X"9"), 42 => Pixel_t'(X"8",X"a",X"9"), 38|44 => Pixel_t'(X"9",X"a",X"a"), 39|43 => Pixel_t'(X"a",X"b",X"b"), 41 => Pixel_t'(X"d",X"e",X"e"), 40 => Pixel_t'(X"f",X"f",X"f")),
    -- 11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|30|31|32|33|34|35|46|47|48|49|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 25|54 => Pixel_t'(X"1",X"1",X"1"), 45 => Pixel_t'(X"1",X"2",X"2"), 29|57 => Pixel_t'(X"2",X"2",X"2"), 26|55 => Pixel_t'(X"3",X"3",X"3"), 27|28|56 => Pixel_t'(X"5",X"5",X"5"), 36|44 => Pixel_t'(X"7",X"7",X"7"), 42 => Pixel_t'(X"8",X"9",X"9"), 38 => Pixel_t'(X"9",X"9",X"9"), 37|39|43 => Pixel_t'(X"9",X"a",X"a"), 40|41 => Pixel_t'(X"e",X"e",X"e")),
    -- 12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|31|32|33|34|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 26|44 => Pixel_t'(X"1",X"1",X"1"), 27|30|35 => Pixel_t'(X"3",X"3",X"3"), 28 => Pixel_t'(X"4",X"5",X"5"), 29 => Pixel_t'(X"5",X"5",X"5"), 36 => Pixel_t'(X"7",X"7",X"7"), 42 => Pixel_t'(X"7",X"8",X"8"), 37|38|39 => Pixel_t'(X"8",X"9",X"9"), 43 => Pixel_t'(X"9",X"9",X"9"), 40 => Pixel_t'(X"9",X"9",X"a"), 41 => Pixel_t'(X"9",X"a",X"a")),
    -- 13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 32 => Pixel_t'(X"0",X"1",X"1"), 33|44 => Pixel_t'(X"1",X"1",X"1"), 28 => Pixel_t'(X"2",X"2",X"3"), 31 => Pixel_t'(X"3",X"4",X"4"), 34 => Pixel_t'(X"4",X"4",X"4"), 29 => Pixel_t'(X"4",X"4",X"5"), 30 => Pixel_t'(X"5",X"5",X"5"), 35|36 => Pixel_t'(X"6",X"7",X"7"), 39 => Pixel_t'(X"7",X"7",X"7"), 37 => Pixel_t'(X"7",X"7",X"8"), 38|40|41|43 => Pixel_t'(X"7",X"8",X"8"), 42 => Pixel_t'(X"8",X"8",X"8")),
    -- 14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 27 => Pixel_t'(X"1",X"1",X"1"), 28|29 => Pixel_t'(X"2",X"2",X"2"), 30 => Pixel_t'(X"3",X"4",X"4"), 35 => Pixel_t'(X"4",X"6",X"6"), 31 => Pixel_t'(X"5",X"5",X"5"), 32|33|34|36|37|38|39|40 => Pixel_t'(X"5",X"6",X"6"), 41 => Pixel_t'(X"6",X"7",X"7"), 42 => Pixel_t'(X"6",X"7",X"8"), 43 => Pixel_t'(X"7",X"8",X"8")),
    -- 15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 45 => Pixel_t'(X"1",X"2",X"2"), 30 => Pixel_t'(X"3",X"3",X"3"), 29 => Pixel_t'(X"3",X"4",X"4"), 21|22|23|31 => Pixel_t'(X"4",X"4",X"4"), 44 => Pixel_t'(X"4",X"5",X"5"), 24|32 => Pixel_t'(X"5",X"6",X"6"), 25 => Pixel_t'(X"6",X"6",X"6"), 28|43 => Pixel_t'(X"6",X"7",X"7"), 26|33|34|42 => Pixel_t'(X"7",X"8",X"8"), 41 => Pixel_t'(X"7",X"8",X"9"), 27|35|36|40 => Pixel_t'(X"8",X"9",X"9"), 37 => Pixel_t'(X"8",X"9",X"a"), 38 => Pixel_t'(X"9",X"a",X"9"), 39 => Pixel_t'(X"9",X"a",X"a")),
    -- 16 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 20 => Pixel_t'(X"4",X"4",X"4"), 45 => Pixel_t'(X"5",X"6",X"6"), 43 => Pixel_t'(X"6",X"7",X"8"), 44 => Pixel_t'(X"6",X"8",X"9"), 42 => Pixel_t'(X"7",X"8",X"9"), 21|22|23|24|25|26|28|29|41 => Pixel_t'(X"9",X"a",X"a"), 30 => Pixel_t'(X"a",X"a",X"a"), 27|31|32|33|34|35|36|37|38 => Pixel_t'(X"a",X"b",X"b"), 39 => Pixel_t'(X"b",X"c",X"b"), 40 => Pixel_t'(X"b",X"c",X"c")),
    -- 17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 45 => Pixel_t'(X"5",X"7",X"7"), 44 => Pixel_t'(X"7",X"8",X"9"), 20 => Pixel_t'(X"8",X"9",X"9"), 35 => Pixel_t'(X"9",X"9",X"9"), 22|23|24|26|30|32|33|34|36 => Pixel_t'(X"9",X"a",X"a"), 43 => Pixel_t'(X"9",X"a",X"b"), 25|27|28|29|37 => Pixel_t'(X"a",X"a",X"a"), 21|31|38|39 => Pixel_t'(X"a",X"b",X"b"), 40 => Pixel_t'(X"c",X"c",X"c"), 42 => Pixel_t'(X"c",X"c",X"d"), 41 => Pixel_t'(X"d",X"e",X"e")),
    -- 18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 19 => Pixel_t'(X"1",X"2",X"2"), 45 => Pixel_t'(X"5",X"6",X"6"), 20 => Pixel_t'(X"7",X"8",X"8"), 44 => Pixel_t'(X"7",X"9",X"9"), 35 => Pixel_t'(X"8",X"7",X"7"), 22|23|25|26|27|28|29|30|32|33|34|36|37|38|39 => Pixel_t'(X"8",X"8",X"8"), 21|24|31 => Pixel_t'(X"8",X"9",X"9"), 40 => Pixel_t'(X"b",X"a",X"a"), 43 => Pixel_t'(X"c",X"d",X"d"), 41|42 => Pixel_t'(X"f",X"d",X"d")),
    -- 19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 21 => Pixel_t'(X"2",X"2",X"2"), 22 => Pixel_t'(X"3",X"3",X"3"), 45 => Pixel_t'(X"4",X"4",X"5"), 23 => Pixel_t'(X"4",X"5",X"5"), 44 => Pixel_t'(X"5",X"6",X"6"), 24 => Pixel_t'(X"6",X"6",X"6"), 27 => Pixel_t'(X"6",X"7",X"6"), 25|26|28|29|30|31|43 => Pixel_t'(X"6",X"7",X"7"), 32|33|34|35 => Pixel_t'(X"7",X"7",X"7"), 36|37 => Pixel_t'(X"7",X"8",X"8"), 38|39 => Pixel_t'(X"8",X"8",X"8"), 40 => Pixel_t'(X"9",X"9",X"9"), 42 => Pixel_t'(X"a",X"9",X"9"), 41 => Pixel_t'(X"b",X"b",X"b")),
    -- 20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 25 => Pixel_t'(X"1",X"2",X"1"), 45 => Pixel_t'(X"2",X"3",X"3"), 26 => Pixel_t'(X"3",X"3",X"3"), 27|28|44 => Pixel_t'(X"3",X"4",X"4"), 29|43 => Pixel_t'(X"4",X"4",X"4"), 30|31 => Pixel_t'(X"4",X"5",X"5"), 42 => Pixel_t'(X"4",X"5",X"6"), 32|33 => Pixel_t'(X"5",X"5",X"5"), 34|35|36 => Pixel_t'(X"5",X"6",X"6"), 41 => Pixel_t'(X"6",X"6",X"6"), 38 => Pixel_t'(X"6",X"6",X"8"), 37|39 => Pixel_t'(X"6",X"7",X"8"), 40 => Pixel_t'(X"7",X"7",X"7")),
    -- 21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 27|28|45 => Pixel_t'(X"1",X"1",X"1"), 29|30|31 => Pixel_t'(X"2",X"2",X"2"), 32 => Pixel_t'(X"2",X"3",X"3"), 33 => Pixel_t'(X"3",X"3",X"3"), 34 => Pixel_t'(X"3",X"3",X"4"), 35|44 => Pixel_t'(X"3",X"4",X"4"), 36|42 => Pixel_t'(X"4",X"4",X"4"), 43 => Pixel_t'(X"4",X"4",X"5"), 41 => Pixel_t'(X"4",X"5",X"5"), 37|38 => Pixel_t'(X"4",X"5",X"6"), 39 => Pixel_t'(X"5",X"5",X"7"), 40 => Pixel_t'(X"5",X"6",X"6")),
    -- 22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 32|33|34|44 => Pixel_t'(X"1",X"1",X"1"), 35 => Pixel_t'(X"2",X"2",X"2"), 36 => Pixel_t'(X"2",X"3",X"3"), 37|41|42 => Pixel_t'(X"3",X"3",X"3"), 38 => Pixel_t'(X"3",X"4",X"3"), 39|40|43 => Pixel_t'(X"4",X"4",X"4")),
    -- 23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 40 => Pixel_t'(X"1",X"1",X"0"), 39 => Pixel_t'(X"1",X"1",X"1"), 37|38 => Pixel_t'(X"2",X"2",X"2")),
    -- 24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")));



    constant pepe_bit_map : bit_map_t (0 to pepe_sizeY-1, 0 to pepe_sizeX-1) :=

    (0 => (48|60 => Pixel_t'("00","01","00"), 27|61|75 => Pixel_t'("01","01","00"), 26|49|59|76 => Pixel_t'("01","01","01"), 28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|62|63|64|65|66|67|68|69|70|71|72|73|74 => Pixel_t'("01","10","01"), 25 => Pixel_t'("10","10","11"), 50|77 => Pixel_t'("10","11","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|51|52|53|54|55|56|57|58|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
1 => (25|58 => Pixel_t'("00","01","00"), 77 => Pixel_t'("00","01","01"), 59 => Pixel_t'("01","01","00"), 26|49|50|76 => Pixel_t'("01","01","01"), 27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75 => Pixel_t'("01","10","01"), 57 => Pixel_t'("01","10","10"), 24|51 => Pixel_t'("10","10","10"), 78 => Pixel_t'("10","10","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|52|53|54|55|56|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
2 => (24|51 => Pixel_t'("00","01","00"), 52|56|57|77|78 => Pixel_t'("01","01","01"), 25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76 => Pixel_t'("01","10","01"), 23|55 => Pixel_t'("10","10","10"), 79 => Pixel_t'("10","11","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|53|54|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
3 => (23|55 => Pixel_t'("00","01","00"), 52 => Pixel_t'("01","01","00"), 53|54|78|79 => Pixel_t'("01","01","01"), 24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77 => Pixel_t'("01","10","01"), 22 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
4 => (22|53|54 => Pixel_t'("00","01","00"), 79 => Pixel_t'("01","01","00"), 23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78 => Pixel_t'("01","10","01"), 80 => Pixel_t'("01","10","10"), 21 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
5 => (21|54|80 => Pixel_t'("00","01","00"), 22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'("01","10","01"), 20|81 => Pixel_t'("10","11","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
6 => (55 => Pixel_t'("01","01","00"), 20|21|54|80 => Pixel_t'("01","01","01"), 81 => Pixel_t'("01","01","10"), 22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'("01","10","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
7 => (55 => Pixel_t'("00","01","00"), 20 => Pixel_t'("01","01","00"), 19|81 => Pixel_t'("01","01","01"), 21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
8 => (39|40|41|42 => Pixel_t'("00","01","00"), 19|38|43|56 => Pixel_t'("01","01","00"), 37|44|45|55|81 => Pixel_t'("01","01","01"), 20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|46|47|48|49|50|51|52|53|54|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 18|82 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
9 => (35|36|45|46|47|56 => Pixel_t'("00","01","00"), 37|44 => Pixel_t'("01","01","00"), 18|34|38|39|40|41|42|43|48|81|82 => Pixel_t'("01","01","01"), 19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|49|50|51|52|53|54|55|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
10 => (33|49|50|56 => Pixel_t'("00","01","00"), 18|32|34|48 => Pixel_t'("01","01","00"), 82 => Pixel_t'("01","01","01"), 19|20|21|22|23|24|25|26|27|28|29|30|31|35|36|37|38|39|40|41|42|43|44|45|46|47|51|52|53|54|55|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81 => Pixel_t'("01","10","01"), 17 => Pixel_t'("01","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
11 => (17|31|51|52 => Pixel_t'("00","01","00"), 32 => Pixel_t'("01","01","00"), 30|50|56|57|82 => Pixel_t'("01","01","01"), 18|19|20|21|22|23|24|25|26|27|28|29|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|53|54|55|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81 => Pixel_t'("01","10","01"), 83 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
12 => (29|30|53|65|66|67|68|69|70|71|72|73|74|75 => Pixel_t'("00","01","00"), 52|57|64|76 => Pixel_t'("01","01","00"), 16|17|54|63|82 => Pixel_t'("01","01","01"), 18|19|20|21|22|23|24|25|26|27|28|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|55|56|58|59|60|61|62|77|78|79|80|81 => Pixel_t'("01","10","01"), 83 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
13 => (28|54|55|57|59|60|61|62|77|78|79|80 => Pixel_t'("00","01","00"), 16|63|76 => Pixel_t'("01","01","00"), 27|29|56|58|64|65|66|75|81|82|83 => Pixel_t'("01","01","01"), 17|18|19|20|21|22|23|24|25|26|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|67|68|69|70|71|72|73|74 => Pixel_t'("01","10","01"), 15 => Pixel_t'("10","11","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
14 => (56|57 => Pixel_t'("00","00","00"), 27|82|84 => Pixel_t'("00","01","00"), 81|83 => Pixel_t'("01","01","00"), 15|16|55|58|59|85 => Pixel_t'("01","01","01"), 17|18|19|20|21|22|23|24|25|26|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 86 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
15 => (57 => Pixel_t'("00","01","00"), 15|86 => Pixel_t'("01","01","00"), 85|87 => Pixel_t'("01","01","01"), 16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84 => Pixel_t'("01","10","01"), 88 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
16 => (58|88 => Pixel_t'("00","01","00"), 15 => Pixel_t'("01","01","00"), 57|87|89 => Pixel_t'("01","01","01"), 16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("01","10","01"), 14 => Pixel_t'("01","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
17 => (59 => Pixel_t'("00","01","00"), 14|58|89|90 => Pixel_t'("01","01","01"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88 => Pixel_t'("01","10","01"), 91 => Pixel_t'("10","10","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
18 => (47|48|49|50|51|52|53|54|55|56|60 => Pixel_t'("00","01","00"), 14|57 => Pixel_t'("01","01","00"), 45|46|58|59|90|91 => Pixel_t'("01","01","01"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("01","10","01"), 13 => Pixel_t'("10","10","10"), 92 => Pixel_t'("10","10","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
19 => (60 => Pixel_t'("00","00","00"), 43|44|45|59|61|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("00","01","00"), 92 => Pixel_t'("00","01","01"), 42|46|58|74|87 => Pixel_t'("01","01","00"), 13|14|47|56|57|62|73|88|91 => Pixel_t'("01","01","01"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|48|49|50|51|52|53|54|55|63|64|65|66|67|68|69|70|71|72|89|90 => Pixel_t'("01","10","01"), 93 => Pixel_t'("10","10","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
20 => (40|41|62|71|72|73|88|89|90|92 => Pixel_t'("00","01","00"), 42|74|87 => Pixel_t'("01","01","00"), 13|39|61|63|70|75|86|91 => Pixel_t'("01","01","01"), 14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|64|65|66|67|68|69|76|77|78|79|80|81|82|83|84|85 => Pixel_t'("01","10","01"), 93 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
21 => (38|39|47|48|49|50|51|52|53|54|55|63|68|69|93 => Pixel_t'("00","01","00"), 13|46|56|70|81|82|92 => Pixel_t'("01","01","00"), 40|45|57|64|67|71|77|78|79|80|83|84|85|91 => Pixel_t'("01","01","01"), 14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|41|42|43|44|58|59|60|61|62|65|66|72|73|74|75|76|86|87|88|89|90 => Pixel_t'("01","10","01"), 94 => Pixel_t'("01","10","10"), 12 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|10|11|95|96|97|98|99 => Pixel_t'("11","11","11")),
22 => (37|43|44|45|58|59|64|66|67|74|75|76|77|85|86|87|88 => Pixel_t'("00","01","00"), 56|57|60|73|78|79|80|81|82|83|84|89 => Pixel_t'("01","01","00"), 12|13|36|38|42|46|55|65|68|72|90|94|95 => Pixel_t'("01","01","01"), 14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|39|40|41|47|48|49|50|51|52|53|54|61|62|63|69|70|71|91|92|93 => Pixel_t'("01","10","01"), 0|1|2|3|4|5|6|7|8|9|10|11|96|97|98|99 => Pixel_t'("11","11","11")),
23 => (12 => Pixel_t'("00","00","00"), 36|41|42|61|62|64|65|70|71|72|90|91 => Pixel_t'("00","01","00"), 35|50|51|52|53|60|69|73|89|92 => Pixel_t'("01","01","00"), 11|40|43|47|48|49|63|74|95|96 => Pixel_t'("01","01","01"), 13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|37|38|39|44|45|46|54|55|56|57|58|59|66|67|68|75|76|77|78|79|80|81|82|83|84|85|86|87|88|93|94 => Pixel_t'("01","10","01"), 10 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|8|9|97|98|99 => Pixel_t'("11","11","11")),
24 => (12|34|40|63|67|68|93|94 => Pixel_t'("00","01","00"), 10|35|39|57|64|66|69|86|88 => Pixel_t'("01","01","00"), 9|11|33|41|43|44|45|46|56|62|70|77|78|79|80|81|82|83|84|85|87|92|95|96 => Pixel_t'("01","01","01"), 13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|36|37|38|42|58|59|60|61|65|71|72|73|74|75|76|89|90|91 => Pixel_t'("01","10","01"), 55 => Pixel_t'("10","10","01"), 8|47|52|53|54 => Pixel_t'("10","10","10"), 0|1|2|3|4|5|6|7|48|49|50|51|97|98|99 => Pixel_t'("11","11","11")),
25 => (79|80|81|82|83 => Pixel_t'("00","00","00"), 8|32|33|38|95 => Pixel_t'("00","01","00"), 48 => Pixel_t'("01","00","01"), 12|31|39|42|60|65|66|74|90 => Pixel_t'("01","01","00"), 37|41|46|47|49|50|58|59|61|75|76|77|78|84|89|94|96 => Pixel_t'("01","01","01"), 9|10|11|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|34|35|36|40|62|63|64|67|68|69|70|71|72|73|88|91|92|93 => Pixel_t'("01","10","01"), 7|43|44|45|57|85|87 => Pixel_t'("10","10","10"), 51 => Pixel_t'("10","10","11"), 0|1|2|3|4|5|6|52|53|54|55|56|86|97|98|99 => Pixel_t'("11","11","11")),
26 => (44|45|46|47|48|49|50|51|77|78|80|81|82|83|84|85 => Pixel_t'("00","00","00"), 7|29|30|37|92|96 => Pixel_t'("00","01","00"), 12|28|31|36|62|63|72 => Pixel_t'("01","01","00"), 11|38|39|40|52|64|73|79|91|97 => Pixel_t'("01","01","01"), 8|9|10|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|32|33|34|35|61|65|66|67|68|69|70|71|93|94|95 => Pixel_t'("01","10","01"), 6|41|43|74|76 => Pixel_t'("10","10","10"), 60 => Pixel_t'("10","11","10"), 0|1|2|3|4|5|42|53|54|55|56|57|58|59|75|86|87|88|89|90|98|99 => Pixel_t'("11","11","11")),
27 => (43|44|47|48|49|50|51|52|76|77|80|81|82|83|84|85|86 => Pixel_t'("00","00","00"), 6|35|65|93 => Pixel_t'("00","01","00"), 34|70|94 => Pixel_t'("01","01","00"), 11|12|36|37|38|64|92|95|97|98 => Pixel_t'("01","01","01"), 7|8|9|10|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|66|67|68|69|71|96 => Pixel_t'("01","10","01"), 5|39|42|53|63|72|75|78 => Pixel_t'("10","10","10"), 0|1|2|3|4|40|41|45|46|54|55|56|57|58|59|60|61|62|73|74|79|87|88|89|90|91|99 => Pixel_t'("11","11","11")),
28 => (42|43|44|47|48|49|50|51|52|53|75|76|77|80|81|82|84|85|86 => Pixel_t'("00","00","00"), 33 => Pixel_t'("00","01","00"), 78 => Pixel_t'("01","00","01"), 11|32|34|66|96 => Pixel_t'("01","01","00"), 5|6|31|36|37|69|79|83|97|98 => Pixel_t'("01","01","01"), 7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|35|67|68|95 => Pixel_t'("01","10","01"), 45|46|65|70|87|94 => Pixel_t'("10","10","10"), 0|1|2|3|4|38|39|40|41|54|55|56|57|58|59|60|61|62|63|64|71|72|73|74|88|89|90|91|92|93|99 => Pixel_t'("11","11","11")),
29 => (42|43|44|45|46|47|48|51|52|53|75|76|77|78|79|80|81|85|86 => Pixel_t'("00","00","00"), 11|26|27|28|29|30|31 => Pixel_t'("00","01","00"), 5|25 => Pixel_t'("01","01","00"), 32|35|66|67|68|84|87|97|98 => Pixel_t'("01","01","01"), 6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24|33|34 => Pixel_t'("01","10","01"), 36 => Pixel_t'("10","10","01"), 4|41|54 => Pixel_t'("10","10","10"), 0|1|2|3|37|38|39|40|49|50|55|56|57|58|59|60|61|62|63|64|65|69|70|71|72|73|74|82|83|88|89|90|91|92|93|94|95|96|99 => Pixel_t'("11","11","11")),
30 => (42|43|44|45|46|47|48|52|53|75|76|77|78|79|80|81|85|86|87 => Pixel_t'("00","00","00"), 11|25 => Pixel_t'("00","01","00"), 67 => Pixel_t'("01","01","00"), 4|34|51|54|66|84|98 => Pixel_t'("01","01","01"), 5|6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24|26|27|28|29|30|31|32|33 => Pixel_t'("01","10","01"), 35|41|74|97 => Pixel_t'("10","10","10"), 0|1|2|3|36|37|38|39|40|49|50|55|56|57|58|59|60|61|62|63|64|65|68|69|70|71|72|73|82|83|88|89|90|91|92|93|94|95|96|99 => Pixel_t'("11","11","11")),
31 => (42|43|44|47|48|51|52|53|54|75|76|77|80|81|82|84|85|86|87 => Pixel_t'("00","00","00"), 78 => Pixel_t'("00","00","01"), 11|25 => Pixel_t'("00","01","00"), 4 => Pixel_t'("01","01","00"), 33|41|45|49|66|83|98 => Pixel_t'("01","01","01"), 46|50 => Pixel_t'("01","01","10"), 5|6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24|26|27|28|29|30|31|32 => Pixel_t'("01","10","01"), 3|34|74 => Pixel_t'("10","10","10"), 79|99 => Pixel_t'("10","10","11"), 0|1|2|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|65|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95|96|97 => Pixel_t'("11","11","11")),
32 => (42|43|44|47|48|49|50|51|52|53|54|75|76|77|78|80|81|82|83|84|85|86|87 => Pixel_t'("00","00","00"), 11|26|27|28 => Pixel_t'("00","01","00"), 29 => Pixel_t'("01","01","00"), 3|25|30|31|32|41|45|79 => Pixel_t'("01","01","01"), 4|5|6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 33|46|66|74|98|99 => Pixel_t'("10","10","10"), 0|1|2|34|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|65|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95|96|97 => Pixel_t'("11","11","11")),
33 => (31|42|43|44|45|46|47|48|49|50|51|52|53|54|75|76|77|78|79|80|81|82|83|84|85|86|87 => Pixel_t'("00","00","00"), 3|30 => Pixel_t'("01","01","00"), 27|28|29|32|41|74|98 => Pixel_t'("01","01","01"), 4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26 => Pixel_t'("01","10","01"), 2|66|99 => Pixel_t'("10","10","10"), 0|1|33|34|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|65|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95|96|97 => Pixel_t'("11","11","11")),
34 => (42|43|44|45|46|47|48|49|50|51|52|53|75|76|77|78|79|80|81|82|83|84|85|86|87 => Pixel_t'("00","00","00"), 32 => Pixel_t'("01","01","00"), 2|3|41|54|98 => Pixel_t'("01","01","01"), 4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31 => Pixel_t'("01","10","01"), 33|65|74|97 => Pixel_t'("10","10","10"), 0|1|34|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|66|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95|96|99 => Pixel_t'("11","11","11")),
35 => (42|43|44|45|46|47|48|49|50|51|52|53|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("00","00","00"), 97 => Pixel_t'("00","00","01"), 2 => Pixel_t'("00","01","00"), 33 => Pixel_t'("01","01","00"), 3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|34|65 => Pixel_t'("01","10","01"), 1|41|54|74|87|96 => Pixel_t'("10","10","10"), 98 => Pixel_t'("10","10","11"), 0|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|66|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95|99 => Pixel_t'("11","11","11")),
36 => (42|43|44|45|46|47|48|49|50|51|52|76|77|78|79|80|81|82|83|84|85|96 => Pixel_t'("00","00","00"), 1|2|34|35|53|64|65|75|86|95 => Pixel_t'("01","01","01"), 3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'("01","10","01"), 36|94 => Pixel_t'("10","10","10"), 97 => Pixel_t'("10","10","11"), 0|37|38|39|40|41|54|55|56|57|58|59|60|61|62|63|66|67|68|69|70|71|72|73|74|87|88|89|90|91|92|93|98|99 => Pixel_t'("11","11","11")),
37 => (43|44|45|46|47|48|49|50|51|52|76|77|78|79|80|81|82|83|84 => Pixel_t'("00","00","00"), 63|93 => Pixel_t'("00","01","00"), 36|65|94 => Pixel_t'("01","01","00"), 1|37|64|66|85|92|95|96 => Pixel_t'("01","01","01"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|62 => Pixel_t'("01","10","01"), 42|91 => Pixel_t'("10","10","10"), 97 => Pixel_t'("10","10","11"), 38 => Pixel_t'("10","11","10"), 0|39|40|41|53|54|55|56|57|58|59|60|61|67|68|69|70|71|72|73|74|75|86|87|88|89|90|98|99 => Pixel_t'("11","11","11")),
38 => (44|45|46|47|48|49|50|78|79|80|81|82|83 => Pixel_t'("00","00","00"), 66|90 => Pixel_t'("00","01","00"), 1|32|38|67|91 => Pixel_t'("01","01","00"), 33|37|39|43|51|61|62|65|68|69|77|84|87|88|89|92|95|96 => Pixel_t'("01","01","01"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|34|35|36|60|63|64|86|93|94 => Pixel_t'("01","10","01"), 70 => Pixel_t'("10","10","01"), 0|40|59|71|85 => Pixel_t'("10","10","10"), 41|42|52|53|54|55|56|57|58|72|73|74|75|76|97|98|99 => Pixel_t'("11","11","11")),
39 => (79|82 => Pixel_t'("00","00","00"), 33|34|65|81|83|94 => Pixel_t'("00","01","00"), 40|58|59|70|71|72|80|84|85|86 => Pixel_t'("01","01","00"), 0|39|41|46|47|57|60|69|73|74|75|78|87|93|95 => Pixel_t'("01","01","01"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|35|36|37|38|61|62|63|64|66|67|68|88|89|90|91|92 => Pixel_t'("01","10","01"), 42|45|48|49|56|76|77 => Pixel_t'("10","10","10"), 43|44|50|51|52|53|54|55|96|97|98|99 => Pixel_t'("11","11","11")),
40 => (0|35|36|64 => Pixel_t'("00","01","00"), 42|43|44|54|55|56 => Pixel_t'("01","01","00"), 34|45|46|47|48|49|50|51|52|53|57|65|78|79|92|93 => Pixel_t'("01","01","01"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|37|38|39|40|41|58|59|60|61|62|63|66|67|68|69|70|71|72|73|74|75|76|77|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 94 => Pixel_t'("10","10","10"), 95|96|97|98|99 => Pixel_t'("11","11","11")),
41 => (37|38|63 => Pixel_t'("00","01","00"), 39 => Pixel_t'("01","01","00"), 0|36|47|48|49|50|51|62|64|92 => Pixel_t'("01","01","01"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|40|41|42|43|44|45|46|52|53|54|55|56|57|58|59|60|61|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
42 => (39|40|41|59|60|61|62 => Pixel_t'("00","01","00"), 42 => Pixel_t'("01","01","00"), 38|58|91 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90 => Pixel_t'("01","10","01"), 92 => Pixel_t'("01","10","10"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
43 => (43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58 => Pixel_t'("00","01","00"), 42 => Pixel_t'("01","01","00"), 41|59|90|91 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("01","10","01"), 92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
44 => (89|90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88 => Pixel_t'("01","10","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
45 => (58 => Pixel_t'("00","01","00"), 57|88 => Pixel_t'("01","01","00"), 89 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87 => Pixel_t'("01","10","01"), 90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
46 => (55 => Pixel_t'("00","01","00"), 56|68|69 => Pixel_t'("01","01","00"), 57|85|86 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|58|59|60|61|62|63|64|65|66|67|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84 => Pixel_t'("01","10","01"), 87 => Pixel_t'("10","10","10"), 88 => Pixel_t'("10","10","11"), 89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
47 => (85 => Pixel_t'("00","00","00"), 54|70|83|84 => Pixel_t'("00","01","00"), 53|55|69|71|82 => Pixel_t'("01","01","00"), 81 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|56|57|58|59|60|61|62|63|64|65|66|67|68|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 86 => Pixel_t'("10","10","10"), 87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
48 => (51|52|72|73|74|75|76|77|78|79|80 => Pixel_t'("00","01","00"), 71|81|82 => Pixel_t'("01","01","00"), 50|53|85|86 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|83|84 => Pixel_t'("01","10","01"), 87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
49 => (74 => Pixel_t'("00","00","00"), 49|50 => Pixel_t'("00","01","00"), 75|86 => Pixel_t'("01","01","00"), 48|51|73|87 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|76|77|78|79|80|81|82|83|84|85 => Pixel_t'("01","10","01"), 88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
50 => (46|47|75 => Pixel_t'("00","01","00"), 48|87 => Pixel_t'("01","01","00"), 49 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("01","10","01"), 88 => Pixel_t'("01","10","10"), 89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
51 => (88 => Pixel_t'("00","01","00"), 46 => Pixel_t'("01","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87 => Pixel_t'("01","10","01"), 89 => Pixel_t'("10","10","10"), 90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
52 => (89 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88 => Pixel_t'("01","10","01"), 90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
53 => (89|90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88 => Pixel_t'("01","10","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
54 => (90 => Pixel_t'("00","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("01","10","01"), 91 => Pixel_t'("10","10","11"), 92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
55 => (90|91 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("01","10","01"), 92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
56 => (91 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90 => Pixel_t'("01","10","01"), 92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
57 => (91 => Pixel_t'("01","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90 => Pixel_t'("01","10","01"), 92 => Pixel_t'("10","10","10"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
58 => (91 => Pixel_t'("01","01","01"), 92 => Pixel_t'("01","01","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90 => Pixel_t'("01","10","01"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
59 => (92 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
60 => (92 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
61 => (92 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
62 => (33|34|35 => Pixel_t'("01","00","00"), 31|32|36|37|38|92 => Pixel_t'("01","01","00"), 30|39|40 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91 => Pixel_t'("01","10","01"), 93 => Pixel_t'("10","10","10"), 94|95|96|97|98|99 => Pixel_t'("11","11","11")),
63 => (30|40|41|92|93 => Pixel_t'("01","00","00"), 29|38|39|42|43|91 => Pixel_t'("01","01","00"), 28|44|45|90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("01","10","01"), 31|32|37 => Pixel_t'("10","01","00"), 33|34|35|36 => Pixel_t'("10","01","01"), 94 => Pixel_t'("10","01","10"), 95|96|97|98|99 => Pixel_t'("11","11","11")),
64 => (28|45|46|90 => Pixel_t'("01","00","00"), 44|47|48|89|94 => Pixel_t'("01","01","00"), 27|49|50|88 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87 => Pixel_t'("01","10","01"), 43|91 => Pixel_t'("10","01","00"), 29|30|31|32|33|34|35|36|37|38|39|40|41|42|92|93 => Pixel_t'("10","01","01"), 95|96|97|98|99 => Pixel_t'("11","11","11")),
65 => (27|49|50|51|87|88 => Pixel_t'("01","00","00"), 48|52|53|86|94 => Pixel_t'("01","01","00"), 26|54|55|85 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84 => Pixel_t'("01","10","01"), 47|89 => Pixel_t'("10","01","00"), 28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|90|91|92|93 => Pixel_t'("10","01","01"), 95 => Pixel_t'("10","10","10"), 96|97|98|99 => Pixel_t'("11","11","11")),
66 => (55|56|84|85 => Pixel_t'("01","00","00"), 26|53|54|57|58|83|94 => Pixel_t'("01","01","00"), 59|60|61|81|82 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'("01","10","01"), 27|30|44|52|86|91 => Pixel_t'("10","01","00"), 28|29|31|32|33|34|35|36|37|38|39|40|41|42|43|45|46|47|48|49|50|51|87|88|89|90|92|93 => Pixel_t'("10","01","01"), 95 => Pixel_t'("10","10","10"), 96|97|98|99 => Pixel_t'("11","11","11")),
67 => (26|61|62|63|80|81 => Pixel_t'("01","00","00"), 59|60|64|65|66|78|79|82 => Pixel_t'("01","01","00"), 25|67|68|69|70|71|72|73|74|75|76|77|94 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 43|44|47|48|49|50|57|58|83|91 => Pixel_t'("10","01","00"), 27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|45|46|51|52|53|54|55|56|84|85|86|87|88|89|90|92|93 => Pixel_t'("10","01","01"), 95|96|97|98|99 => Pixel_t'("11","11","11")),
68 => (32|33|34|35|36|37|38|39|70|71|72|74|75|93 => Pixel_t'("01","00","00"), 25|66|67|68|69|73|76|77 => Pixel_t'("01","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 26|31|50|51|52|53|54|56|57|63|64|65|78|79 => Pixel_t'("10","01","00"), 27|28|29|30|40|41|42|43|44|45|46|47|48|49|55|58|59|60|61|62|80|81|82|83|84|85|86|87|88|89|90|91|92 => Pixel_t'("10","01","01"), 94 => Pixel_t'("10","10","10"), 95|96|97|98|99 => Pixel_t'("11","11","11")),
69 => (40|41|42|43|92 => Pixel_t'("01","00","00"), 25|44 => Pixel_t'("01","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 38|39|54|59|62|79|80|81|88 => Pixel_t'("10","01","00"), 26|27|28|29|30|31|32|33|34|35|36|37|45|46|47|48|49|50|51|52|53|55|56|57|58|60|61|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|82|83|84|85|86|87|89|90|91 => Pixel_t'("10","01","01"), 93 => Pixel_t'("10","10","10"), 94|95|96|97|98|99 => Pixel_t'("11","11","11")),
70 => (44|45|46|47|48 => Pixel_t'("01","00","00"), 25 => Pixel_t'("01","01","00"), 90|91 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 32|43|49|78|79 => Pixel_t'("10","01","00"), 26|27|28|29|30|31|33|34|35|36|37|38|39|40|41|42|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|80|81|82|83|84|85|86|87|88|89 => Pixel_t'("10","01","01"), 92 => Pixel_t'("10","10","10"), 93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
71 => (49|50|51|52|53|89 => Pixel_t'("01","00","00"), 25|54|87|88 => Pixel_t'("01","01","00"), 90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 29|48 => Pixel_t'("10","01","00"), 26|27|28|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("10","01","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
72 => (55|56|57|58|59|60|81|82|83|84|85|86 => Pixel_t'("01","00","00"), 25|26|54|61|62|63|78|79|80|87|89 => Pixel_t'("01","01","00"), 90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'("01","10","01"), 42|43|44|52|53|64|65|66|76|77|88 => Pixel_t'("10","01","00"), 27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|45|46|47|48|49|50|51|67|68|69|70|71|72|73|74|75 => Pixel_t'("10","01","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
73 => (65|66|67|68|69|70|71|72|73|74|75|76 => Pixel_t'("01","00","00"), 26|64|77|78|90 => Pixel_t'("01","01","00"), 27 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25 => Pixel_t'("01","10","01"), 44|45|59|60|61|62|63|79|80|81 => Pixel_t'("10","01","00"), 28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|46|47|48|49|50|51|52|53|54|55|56|57|58|82|83|84|85|86|87|88|89 => Pixel_t'("10","01","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
74 => (28 => Pixel_t'("00","00","00"), 21|27 => Pixel_t'("00","01","00"), 32|33|34|35|36 => Pixel_t'("01","00","00"), 29|30|31|37|38|39|90 => Pixel_t'("01","01","00"), 40 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|22|23|24|25|26 => Pixel_t'("01","10","01"), 47|48|49|85|86|87 => Pixel_t'("10","01","00"), 41|42|43|44|45|46|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|88|89 => Pixel_t'("10","01","01"), 91 => Pixel_t'("10","10","10"), 92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
75 => (21|39|40|41|42|43|44 => Pixel_t'("01","01","00"), 22|37|38|90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|23|24|25|26|27|28|29|30|31|32|33|34|35|36 => Pixel_t'("01","10","01"), 59|60|83|87 => Pixel_t'("10","01","00"), 45|46|47|48|49|50|51|52|53|54|55|56|57|58|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|84|85|86|88|89 => Pixel_t'("10","01","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
76 => (22 => Pixel_t'("00","01","00"), 44|45|46|47|48 => Pixel_t'("01","01","00"), 43|49|89|90 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42 => Pixel_t'("01","10","01"), 59|60|61|63|71|86|87 => Pixel_t'("10","01","00"), 50|51|52|53|54|55|56|57|58|62|64|65|66|67|68|69|70|72|73|74|75|76|77|78|79|80|81|82|83|84|85|88 => Pixel_t'("10","01","01"), 91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
77 => (50 => Pixel_t'("00","01","00"), 22|23|48|49|51|52|53 => Pixel_t'("01","01","00"), 47|54|88|89 => Pixel_t'("01","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46 => Pixel_t'("01","10","01"), 74|75|76|77|78|79|82 => Pixel_t'("10","01","00"), 55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|80|81|83|84|85|86|87 => Pixel_t'("10","01","01"), 90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
78 => (23|24|55|56 => Pixel_t'("00","01","00"), 53|54|57|58|59|60|61|62|63|87 => Pixel_t'("01","01","00"), 0|52|64|88 => Pixel_t'("01","01","01"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51 => Pixel_t'("01","10","01"), 65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'("10","01","01"), 89 => Pixel_t'("10","10","11"), 90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
79 => (25|65|66|67|68|69|70|71 => Pixel_t'("00","01","00"), 83 => Pixel_t'("01","00","00"), 24|26|60|61|62|63|64|72|73|74|75|76|77|78|79|80|81|82 => Pixel_t'("01","01","00"), 1|27|59|84|85|86 => Pixel_t'("01","01","01"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58 => Pixel_t'("01","10","01"), 0|87 => Pixel_t'("10","10","10"), 88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
80 => (81 => Pixel_t'("00","00","00"), 27 => Pixel_t'("00","01","00"), 26|28 => Pixel_t'("01","01","00"), 1|2|74|75|76|77|78|79|80|82 => Pixel_t'("01","01","01"), 3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("01","10","01"), 83|84 => Pixel_t'("10","10","11"), 0|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
81 => (2 => Pixel_t'("00","00","00"), 3|80 => Pixel_t'("01","01","01"), 81 => Pixel_t'("01","01","10"), 4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'("01","10","01"), 1 => Pixel_t'("10","10","10"), 0|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
82 => (1 => Pixel_t'("00","00","01"), 4 => Pixel_t'("00","01","00"), 3|79 => Pixel_t'("01","01","00"), 2|5 => Pixel_t'("01","01","01"), 0 => Pixel_t'("01","01","10"), 6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78 => Pixel_t'("01","10","01"), 80 => Pixel_t'("01","10","10"), 81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
83 => (2 => Pixel_t'("00","00","01"), 1 => Pixel_t'("00","00","10"), 0 => Pixel_t'("00","00","11"), 5|6|78 => Pixel_t'("00","01","00"), 3|4|77 => Pixel_t'("01","01","01"), 7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76 => Pixel_t'("01","10","01"), 79 => Pixel_t'("10","10","10"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
84 => (3 => Pixel_t'("00","00","01"), 7|8 => Pixel_t'("00","01","00"), 0|1|2 => Pixel_t'("00","01","11"), 4|6|9|76|77 => Pixel_t'("01","01","01"), 5|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75 => Pixel_t'("01","10","01"), 78 => Pixel_t'("10","10","10"), 79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
85 => (4 => Pixel_t'("00","00","10"), 9|10|75 => Pixel_t'("00","01","00"), 5 => Pixel_t'("00","01","01"), 0|1|2|3 => Pixel_t'("00","01","11"), 8|11|74|76 => Pixel_t'("01","01","01"), 6|7|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("01","10","01"), 77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
86 => (6 => Pixel_t'("00","00","01"), 5 => Pixel_t'("00","00","11"), 12|13 => Pixel_t'("00","01","00"), 0|1|2|3|4 => Pixel_t'("00","01","11"), 11|73 => Pixel_t'("01","01","00"), 7|10|14|72|74 => Pixel_t'("01","01","01"), 8|9|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71 => Pixel_t'("01","10","01"), 75 => Pixel_t'("10","10","10"), 76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
87 => (8 => Pixel_t'("00","00","01"), 7 => Pixel_t'("00","00","10"), 14|15|16|71 => Pixel_t'("00","01","00"), 0|1|2|3|4|5|6 => Pixel_t'("00","01","11"), 13 => Pixel_t'("01","01","00"), 9|17|70|72 => Pixel_t'("01","01","01"), 10|11|12|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69 => Pixel_t'("01","10","01"), 73 => Pixel_t'("10","10","10"), 74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
88 => (9 => Pixel_t'("00","00","10"), 8 => Pixel_t'("00","00","11"), 17|18|19|20|69 => Pixel_t'("00","01","00"), 10 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7 => Pixel_t'("00","01","11"), 16|21 => Pixel_t'("01","01","00"), 11|22|67|68|70 => Pixel_t'("01","01","01"), 12|13|14|15|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66 => Pixel_t'("01","10","01"), 71 => Pixel_t'("10","10","10"), 72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
89 => (11 => Pixel_t'("00","00","10"), 10 => Pixel_t'("00","00","11"), 22|23|24|25|26 => Pixel_t'("00","01","00"), 12 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7|8|9 => Pixel_t'("00","01","11"), 21|27 => Pixel_t'("01","01","00"), 13|28|29|66|67 => Pixel_t'("01","01","01"), 14|15|16|17|18|19|20|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65 => Pixel_t'("01","10","01"), 68|69 => Pixel_t'("10","10","10"), 70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
90 => (14|64|65 => Pixel_t'("00","00","01"), 13 => Pixel_t'("00","00","10"), 12 => Pixel_t'("00","00","11"), 29|30|31|32|33|63 => Pixel_t'("00","01","00"), 0|1|2|3|4|5|6|7|8|9|10|11 => Pixel_t'("00","01","11"), 27|28|34|35|61|62 => Pixel_t'("01","01","00"), 15|36|37|38|60|66 => Pixel_t'("01","01","01"), 16|17|18|19|20|21|22|23|24|25|26|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59 => Pixel_t'("01","10","01"), 67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
91 => (15|16|64|65 => Pixel_t'("00","00","10"), 37|38|39|40|41|42|43|44|45|46|47|48|50|51|52|53|54|55|56|57|58|59|60 => Pixel_t'("00","01","00"), 17 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","01","11"), 35|36|49|61 => Pixel_t'("01","01","00"), 18|34|62|63 => Pixel_t'("01","01","01"), 66 => Pixel_t'("01","01","10"), 19|20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'("01","10","01"), 67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
92 => (19 => Pixel_t'("00","00","01"), 18|63|66 => Pixel_t'("00","00","10"), 17 => Pixel_t'("00","00","11"), 20 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|64|65 => Pixel_t'("00","01","11"), 21|22|47|48|49|50|51|62 => Pixel_t'("01","01","01"), 67 => Pixel_t'("01","01","10"), 23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|52|53|54|55|56|57|58|59|60|61 => Pixel_t'("01","10","01"), 68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
93 => (23 => Pixel_t'("00","00","01"), 21|22|62|67 => Pixel_t'("00","00","10"), 20|63 => Pixel_t'("00","00","11"), 24|25|61 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|64|65|66 => Pixel_t'("00","01","11"), 26|27|28|60 => Pixel_t'("01","01","01"), 68 => Pixel_t'("01","01","10"), 29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59 => Pixel_t'("01","10","01"), 69 => Pixel_t'("10","10","11"), 70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
94 => (31 => Pixel_t'("00","00","01"), 25|26|27|28|29|30|59|60|69 => Pixel_t'("00","00","10"), 24|61|68 => Pixel_t'("00","00","11"), 32|33|58 => Pixel_t'("00","01","01"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|62|63|64|65|66|67 => Pixel_t'("00","01","11"), 34|35|36|37|38|39|54|55|56|57 => Pixel_t'("01","01","01"), 40|41|42|43|44|45|46|47|48|49|50|51|52|53 => Pixel_t'("01","10","01"), 70 => Pixel_t'("10","10","10"), 71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
95 => (43|44|51 => Pixel_t'("00","00","01"), 34|35|36|37|38|39|40|41|42|52|53|54|55|56|70 => Pixel_t'("00","00","10"), 32|33|57|58 => Pixel_t'("00","00","11"), 45|48|49|50 => Pixel_t'("00","01","01"), 46|47 => Pixel_t'("00","01","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|59|60|61|62|63|64|65|66|67|68|69 => Pixel_t'("00","01","11"), 71 => Pixel_t'("01","01","10"), 72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
96 => (71|72 => Pixel_t'("00","00","10"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70 => Pixel_t'("00","01","11"), 73 => Pixel_t'("10","10","11"), 74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
97 => (73 => Pixel_t'("00","00","10"), 72 => Pixel_t'("00","00","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71 => Pixel_t'("00","01","11"), 74 => Pixel_t'("10","10","11"), 75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
98 => (74 => Pixel_t'("00","00","10"), 73 => Pixel_t'("00","00","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72 => Pixel_t'("00","01","11"), 75 => Pixel_t'("10","10","11"), 76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")),
99 => (75 => Pixel_t'("00","00","10"), 74 => Pixel_t'("00","00","11"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","01","11"), 76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'("11","11","11")));




end package;