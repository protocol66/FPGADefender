(0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
1 => (0|1|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 2|3|4|5 => Pixel_t'("11","11","11")),
2 => (0|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3|4 => Pixel_t'("11","11","11")),
3 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
4 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
5 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
6 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
7 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
8 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
9 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
10 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
11 => (0|4|13|14 => Pixel_t'("00","00","00"), 1|2|3|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
14 => (0|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|4|11|12|13 => Pixel_t'("11","11","11")),
15 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
20 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));