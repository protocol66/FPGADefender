library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.my_data_types.all;

package bitmaps is
    constant BACKGROUND : Pixel_t := BLACK;
    constant MAIN_CLK_FREQ : integer := 50000000;

    constant screen_HEIGHT : positive := 479;
    constant screen_WIDTH : positive := 639;

    constant pepe_sizeX : positive := 100;
    constant pepe_sizeY : positive := 100;

    constant line_sizeX : positive := screen_WIDTH;
    constant line_sizeY : positive := 2;

    constant ship_sizeX : positive := 25;
    constant ship_sizeY : positive := 25;
    
    constant laser_sizeX : positive := ship_sizeX;
    constant laser_sizeY : positive := 1;

    constant score_sizeX : positive := 15;
    constant score_sizeY : positive := 25;
    constant score_space_size :positive := 5;
    constant score_board_sizeX : positive := (score_sizeX + score_space_size)*5 + score_sizeY;
    constant score_board_sizeY : positive := score_sizeY;

    constant alien1_sizeX : positive := 30;
    constant alien1_sizeY : positive := 30;

    constant alien2_sizeX : positive := 20;
    constant alien2_sizeY : positive := 20;

    constant alien3_sizeX : positive := 10;
    constant alien3_sizeY : positive := 10;

    constant asteroid_sizeX : positive := 40;
    constant asteroid_sizeY : positive := 40;

    constant H_LINE : bit_map_t (0 to line_sizeY-1, 0 to line_sizeX-1) := (others => (others => WHITE));
    constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) := (others => (others => TEAL));
    constant LASER : bit_map_t (0 to laser_sizeY-1, 0 to laser_sizeX-1) := (others => (others => GREEN));
    constant ALIEN_1 : bit_map_t (0 to alien1_sizeY-1, 0 to alien1_sizeX-1) := (others => (others => YELLOW));
    constant ALIEN_2 : bit_map_t (0 to alien2_sizeY-1, 0 to alien2_sizeX-1) := (others => (others => RED)); 
    constant ALIEN_3 : bit_map_t (0 to alien3_sizeY-1, 0 to alien3_sizeX-1) := (others => (others => BLUE));  
    constant ASTEROID : bit_map_t (0 to asteroid_sizeY-1, 0 to asteroid_sizeX-1) := (others => (others => PURPLE)); 
    constant SATELLITE : bit_map_t (0 to asteroid_sizeY-1, 0 to asteroid_sizeX-1) := (others => (others => GREEN)); 

    constant fx1 : Sound_FX_t := (18, (550, 404, 315, 494, 182, 260, 455, 387, 340, 550, 404, 315, 494, 182, 260, 455, 387, 340, others => 0));
    constant fx2 : Sound_FX_t := (10, (300, 350, 500, 700, 990, 970, 1050, 1010, 950, 800, 770, 640, 500, 350, 355, others => 0));
    constant fx3 : Sound_FX_t := (6,  (500, 790, 950, 1300, 1710, 1650, 1300, 800, 700, others=> 0));
    constant fx4 : Sound_FX_t := (60, (1300, 1650, 1660, 1510, 1309, 1158, 1007, 855, others=> 0));
    constant fx5 : Sound_FX_t := (25, (300, 210, 310, 170, 250, 210, 310, 120, 220, 170, 160, 90, 290, 230, 140, 320, 200, 100, 250, 290, others => 0));
    constant fx6 : Sound_FX_t := (15, (700, 702, 698, 701, 699, 700, 250, 251, 249, 252, 248, 130, 131, 129, 132, 128, 130, 130, others=>0));

    -- constant score_9 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    -- constant score_8 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    -- constant score_7 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    -- constant score_6 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    -- constant score_5 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => PURPLE));
    -- constant score_4 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => YELLOW));
    -- constant score_3 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    -- constant score_2 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    -- constant score_1 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    -- constant score_0 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    constant score_blank : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BACKGROUND));
    
    -- DONT USE THIS... adds 30+ min to compile time...
    -- constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) :=
    -- (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")),
    -- 1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")),
    -- 2 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 1|2|3|4 => Pixel_t'(X"1",X"1",X"1"), 5|57 => Pixel_t'(X"2",X"2",X"2"), 54 => Pixel_t'(X"3",X"3",X"3"), 55 => Pixel_t'(X"3",X"4",X"4"), 6|36 => Pixel_t'(X"5",X"5",X"6"), 56 => Pixel_t'(X"5",X"6",X"6"), 11|12|13|14|15|31|32|33|34 => Pixel_t'(X"6",X"7",X"7"), 7|8|9|10|16|35 => Pixel_t'(X"7",X"7",X"7"), 19|20|22|24|25 => Pixel_t'(X"7",X"7",X"8"), 17|18|21|23|26|27|28|29|30 => Pixel_t'(X"7",X"8",X"8")),
    -- 3 => (38|39|40|41|42|43|44|45|46|47|48|49|50|51|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 0|37|52 => Pixel_t'(X"1",X"1",X"1"), 58 => Pixel_t'(X"2",X"2",X"2"), 53 => Pixel_t'(X"3",X"3",X"3"), 21|22|23|29 => Pixel_t'(X"6",X"6",X"6"), 19|20|24|25|26|28 => Pixel_t'(X"6",X"6",X"7"), 17|18|27 => Pixel_t'(X"6",X"7",X"7"), 1|16|32 => Pixel_t'(X"7",X"7",X"7"), 15 => Pixel_t'(X"7",X"7",X"8"), 14|30|54 => Pixel_t'(X"7",X"8",X"8"), 2 => Pixel_t'(X"8",X"8",X"8"), 4|5|13|31|33|34|35 => Pixel_t'(X"8",X"8",X"9"), 3|36|55|57 => Pixel_t'(X"8",X"9",X"9"), 12 => Pixel_t'(X"9",X"9",X"a"), 6|56 => Pixel_t'(X"9",X"a",X"a"), 7|8 => Pixel_t'(X"a",X"a",X"b"), 11 => Pixel_t'(X"b",X"b",X"c"), 9 => Pixel_t'(X"b",X"c",X"c"), 10 => Pixel_t'(X"c",X"d",X"d")),
    -- 4 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 20|21|23|26|27|28 => Pixel_t'(X"1",X"1",X"1"), 16|17|18|19|22|24|25 => Pixel_t'(X"1",X"1",X"2"), 12|13|14|15|32|51 => Pixel_t'(X"2",X"2",X"2"), 1|29|59 => Pixel_t'(X"3",X"3",X"3"), 11 => Pixel_t'(X"4",X"4",X"4"), 33 => Pixel_t'(X"5",X"5",X"6"), 31|36|52 => Pixel_t'(X"5",X"6",X"6"), 5 => Pixel_t'(X"6",X"6",X"7"), 2|30 => Pixel_t'(X"6",X"7",X"7"), 55 => Pixel_t'(X"7",X"7",X"7"), 3|4|34|35|53|54|56|58 => Pixel_t'(X"7",X"8",X"8"), 6 => Pixel_t'(X"8",X"8",X"9"), 57 => Pixel_t'(X"8",X"9",X"9"), 7 => Pixel_t'(X"9",X"9",X"9"), 8 => Pixel_t'(X"9",X"a",X"a"), 10 => Pixel_t'(X"a",X"b",X"b"), 9 => Pixel_t'(X"c",X"d",X"d")),
    -- 5 => (0|1|37|38|39|40|41|42|43|44|45|46|47|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 48|63 => Pixel_t'(X"1",X"1",X"1"), 36|49|62 => Pixel_t'(X"2",X"2",X"2"), 21|22|23 => Pixel_t'(X"2",X"3",X"3"), 16|17|18|19|20|24|25|26|27|28 => Pixel_t'(X"3",X"3",X"3"), 15 => Pixel_t'(X"3",X"3",X"4"), 14 => Pixel_t'(X"3",X"4",X"4"), 2|13|32|61 => Pixel_t'(X"4",X"4",X"4"), 12|31 => Pixel_t'(X"4",X"4",X"5"), 50 => Pixel_t'(X"4",X"5",X"5"), 3|11|29 => Pixel_t'(X"5",X"6",X"6"), 30 => Pixel_t'(X"6",X"6",X"6"), 51|60 => Pixel_t'(X"6",X"7",X"7"), 4|5|33|52|55 => Pixel_t'(X"7",X"7",X"7"), 6|10|53|54 => Pixel_t'(X"7",X"7",X"8"), 7|9|34|35|56|59 => Pixel_t'(X"7",X"8",X"8"), 8 => Pixel_t'(X"8",X"8",X"8"), 58 => Pixel_t'(X"8",X"9",X"9"), 57 => Pixel_t'(X"9",X"a",X"a")),
    -- 6 => (0|1|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 2 => Pixel_t'(X"0",X"1",X"0"), 6|7|8|9|72 => Pixel_t'(X"1",X"1",X"1"), 68|69|70|71 => Pixel_t'(X"2",X"2",X"2"), 5 => Pixel_t'(X"2",X"2",X"3"), 10 => Pixel_t'(X"2",X"3",X"3"), 44|67 => Pixel_t'(X"3",X"3",X"3"), 4|45 => Pixel_t'(X"3",X"4",X"4"), 29|30|31|32|66 => Pixel_t'(X"4",X"4",X"4"), 15|16 => Pixel_t'(X"4",X"4",X"5"), 3|11|14|33|34|43|46 => Pixel_t'(X"4",X"5",X"5"), 38 => Pixel_t'(X"4",X"7",X"8"), 12|13|19|20|21|22|23|24|28|35|40 => Pixel_t'(X"5",X"5",X"5"), 25|65 => Pixel_t'(X"5",X"5",X"6"), 17|18|26|27|41|47 => Pixel_t'(X"5",X"6",X"6"), 42 => Pixel_t'(X"5",X"7",X"7"), 39 => Pixel_t'(X"6",X"6",X"6"), 48|51|52|53|54|55|56|57|58|64 => Pixel_t'(X"6",X"7",X"7"), 49|50|59|63 => Pixel_t'(X"7",X"7",X"7"), 60|61|62 => Pixel_t'(X"7",X"8",X"8")),
    -- 7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|29|30|31|32|33|34|35|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 17|28 => Pixel_t'(X"2",X"2",X"2"), 18|19|26|43 => Pixel_t'(X"3",X"3",X"3"), 44 => Pixel_t'(X"3",X"3",X"4"), 25|27|42|45 => Pixel_t'(X"3",X"4",X"4"), 38 => Pixel_t'(X"3",X"6",X"6"), 20 => Pixel_t'(X"4",X"4",X"4"), 46 => Pixel_t'(X"4",X"4",X"5"), 21|22|24|41|47|48|49 => Pixel_t'(X"4",X"5",X"5"), 23 => Pixel_t'(X"5",X"5",X"5"), 53 => Pixel_t'(X"5",X"5",X"6"), 50|51|52|54|55|57 => Pixel_t'(X"5",X"6",X"6"), 56 => Pixel_t'(X"6",X"6",X"6"), 58|72 => Pixel_t'(X"6",X"6",X"7"), 59 => Pixel_t'(X"7",X"7",X"8"), 39|40|60|61|62|68|71 => Pixel_t'(X"7",X"8",X"8"), 69|70 => Pixel_t'(X"8",X"8",X"9"), 63|64|67 => Pixel_t'(X"8",X"9",X"9"), 65|66 => Pixel_t'(X"8",X"9",X"a")),
    -- 8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|27|28|29|30|31|32|33|34|35|36|37|73 => Pixel_t'(X"0",X"0",X"0"), 26 => Pixel_t'(X"0",X"1",X"0"), 20|38 => Pixel_t'(X"1",X"1",X"1"), 50|51|52 => Pixel_t'(X"2",X"2",X"2"), 68 => Pixel_t'(X"2",X"3",X"3"), 21|49|53|64|65|66|67|69|70|71|72 => Pixel_t'(X"3",X"3",X"3"), 63 => Pixel_t'(X"3",X"3",X"4"), 25|59|60 => Pixel_t'(X"3",X"4",X"4"), 22|23|54|57|58|61|62 => Pixel_t'(X"4",X"4",X"4"), 55 => Pixel_t'(X"4",X"5",X"4"), 24|48|56 => Pixel_t'(X"4",X"5",X"5"), 42|45|46|47 => Pixel_t'(X"5",X"6",X"6"), 43|44 => Pixel_t'(X"6",X"6",X"6"), 39 => Pixel_t'(X"6",X"7",X"6"), 40|41 => Pixel_t'(X"7",X"8",X"8")),
    -- 9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|28|29|30|31|32|33|34|35|36|50|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 49 => Pixel_t'(X"0",X"1",X"1"), 21|27|37|48|51|52|53|61 => Pixel_t'(X"1",X"1",X"1"), 22|23 => Pixel_t'(X"2",X"2",X"2"), 58|59|60 => Pixel_t'(X"3",X"3",X"3"), 24 => Pixel_t'(X"3",X"4",X"4"), 26|54 => Pixel_t'(X"4",X"4",X"4"), 25 => Pixel_t'(X"4",X"5",X"5"), 47|57 => Pixel_t'(X"5",X"5",X"5"), 38 => Pixel_t'(X"7",X"8",X"8"), 55|56 => Pixel_t'(X"8",X"8",X"8"), 39|45|46 => Pixel_t'(X"8",X"9",X"9"), 42 => Pixel_t'(X"8",X"a",X"9"), 44 => Pixel_t'(X"9",X"a",X"a"), 43 => Pixel_t'(X"a",X"a",X"a"), 40|41 => Pixel_t'(X"c",X"d",X"d")),
    -- 10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|29|30|31|32|33|34|35|36|47|48|49|50|51|52|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 24|53|59 => Pixel_t'(X"1",X"1",X"1"), 28 => Pixel_t'(X"1",X"2",X"2"), 54 => Pixel_t'(X"2",X"2",X"2"), 25 => Pixel_t'(X"3",X"4",X"4"), 46|57|58 => Pixel_t'(X"4",X"4",X"4"), 27 => Pixel_t'(X"4",X"5",X"5"), 26 => Pixel_t'(X"5",X"5",X"5"), 37|55 => Pixel_t'(X"7",X"8",X"8"), 45 => Pixel_t'(X"8",X"8",X"8"), 56 => Pixel_t'(X"8",X"9",X"9"), 42 => Pixel_t'(X"8",X"a",X"9"), 38|44 => Pixel_t'(X"9",X"a",X"a"), 39|43 => Pixel_t'(X"a",X"b",X"b"), 41 => Pixel_t'(X"d",X"e",X"e"), 40 => Pixel_t'(X"f",X"f",X"f")),
    -- 11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|30|31|32|33|34|35|46|47|48|49|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 25|54 => Pixel_t'(X"1",X"1",X"1"), 45 => Pixel_t'(X"1",X"2",X"2"), 29|57 => Pixel_t'(X"2",X"2",X"2"), 26|55 => Pixel_t'(X"3",X"3",X"3"), 27|28|56 => Pixel_t'(X"5",X"5",X"5"), 36|44 => Pixel_t'(X"7",X"7",X"7"), 42 => Pixel_t'(X"8",X"9",X"9"), 38 => Pixel_t'(X"9",X"9",X"9"), 37|39|43 => Pixel_t'(X"9",X"a",X"a"), 40|41 => Pixel_t'(X"e",X"e",X"e")),
    -- 12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|31|32|33|34|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 26|44 => Pixel_t'(X"1",X"1",X"1"), 27|30|35 => Pixel_t'(X"3",X"3",X"3"), 28 => Pixel_t'(X"4",X"5",X"5"), 29 => Pixel_t'(X"5",X"5",X"5"), 36 => Pixel_t'(X"7",X"7",X"7"), 42 => Pixel_t'(X"7",X"8",X"8"), 37|38|39 => Pixel_t'(X"8",X"9",X"9"), 43 => Pixel_t'(X"9",X"9",X"9"), 40 => Pixel_t'(X"9",X"9",X"a"), 41 => Pixel_t'(X"9",X"a",X"a")),
    -- 13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 32 => Pixel_t'(X"0",X"1",X"1"), 33|44 => Pixel_t'(X"1",X"1",X"1"), 28 => Pixel_t'(X"2",X"2",X"3"), 31 => Pixel_t'(X"3",X"4",X"4"), 34 => Pixel_t'(X"4",X"4",X"4"), 29 => Pixel_t'(X"4",X"4",X"5"), 30 => Pixel_t'(X"5",X"5",X"5"), 35|36 => Pixel_t'(X"6",X"7",X"7"), 39 => Pixel_t'(X"7",X"7",X"7"), 37 => Pixel_t'(X"7",X"7",X"8"), 38|40|41|43 => Pixel_t'(X"7",X"8",X"8"), 42 => Pixel_t'(X"8",X"8",X"8")),
    -- 14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 27 => Pixel_t'(X"1",X"1",X"1"), 28|29 => Pixel_t'(X"2",X"2",X"2"), 30 => Pixel_t'(X"3",X"4",X"4"), 35 => Pixel_t'(X"4",X"6",X"6"), 31 => Pixel_t'(X"5",X"5",X"5"), 32|33|34|36|37|38|39|40 => Pixel_t'(X"5",X"6",X"6"), 41 => Pixel_t'(X"6",X"7",X"7"), 42 => Pixel_t'(X"6",X"7",X"8"), 43 => Pixel_t'(X"7",X"8",X"8")),
    -- 15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 45 => Pixel_t'(X"1",X"2",X"2"), 30 => Pixel_t'(X"3",X"3",X"3"), 29 => Pixel_t'(X"3",X"4",X"4"), 21|22|23|31 => Pixel_t'(X"4",X"4",X"4"), 44 => Pixel_t'(X"4",X"5",X"5"), 24|32 => Pixel_t'(X"5",X"6",X"6"), 25 => Pixel_t'(X"6",X"6",X"6"), 28|43 => Pixel_t'(X"6",X"7",X"7"), 26|33|34|42 => Pixel_t'(X"7",X"8",X"8"), 41 => Pixel_t'(X"7",X"8",X"9"), 27|35|36|40 => Pixel_t'(X"8",X"9",X"9"), 37 => Pixel_t'(X"8",X"9",X"a"), 38 => Pixel_t'(X"9",X"a",X"9"), 39 => Pixel_t'(X"9",X"a",X"a")),
    -- 16 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 20 => Pixel_t'(X"4",X"4",X"4"), 45 => Pixel_t'(X"5",X"6",X"6"), 43 => Pixel_t'(X"6",X"7",X"8"), 44 => Pixel_t'(X"6",X"8",X"9"), 42 => Pixel_t'(X"7",X"8",X"9"), 21|22|23|24|25|26|28|29|41 => Pixel_t'(X"9",X"a",X"a"), 30 => Pixel_t'(X"a",X"a",X"a"), 27|31|32|33|34|35|36|37|38 => Pixel_t'(X"a",X"b",X"b"), 39 => Pixel_t'(X"b",X"c",X"b"), 40 => Pixel_t'(X"b",X"c",X"c")),
    -- 17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 45 => Pixel_t'(X"5",X"7",X"7"), 44 => Pixel_t'(X"7",X"8",X"9"), 20 => Pixel_t'(X"8",X"9",X"9"), 35 => Pixel_t'(X"9",X"9",X"9"), 22|23|24|26|30|32|33|34|36 => Pixel_t'(X"9",X"a",X"a"), 43 => Pixel_t'(X"9",X"a",X"b"), 25|27|28|29|37 => Pixel_t'(X"a",X"a",X"a"), 21|31|38|39 => Pixel_t'(X"a",X"b",X"b"), 40 => Pixel_t'(X"c",X"c",X"c"), 42 => Pixel_t'(X"c",X"c",X"d"), 41 => Pixel_t'(X"d",X"e",X"e")),
    -- 18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 19 => Pixel_t'(X"1",X"2",X"2"), 45 => Pixel_t'(X"5",X"6",X"6"), 20 => Pixel_t'(X"7",X"8",X"8"), 44 => Pixel_t'(X"7",X"9",X"9"), 35 => Pixel_t'(X"8",X"7",X"7"), 22|23|25|26|27|28|29|30|32|33|34|36|37|38|39 => Pixel_t'(X"8",X"8",X"8"), 21|24|31 => Pixel_t'(X"8",X"9",X"9"), 40 => Pixel_t'(X"b",X"a",X"a"), 43 => Pixel_t'(X"c",X"d",X"d"), 41|42 => Pixel_t'(X"f",X"d",X"d")),
    -- 19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 21 => Pixel_t'(X"2",X"2",X"2"), 22 => Pixel_t'(X"3",X"3",X"3"), 45 => Pixel_t'(X"4",X"4",X"5"), 23 => Pixel_t'(X"4",X"5",X"5"), 44 => Pixel_t'(X"5",X"6",X"6"), 24 => Pixel_t'(X"6",X"6",X"6"), 27 => Pixel_t'(X"6",X"7",X"6"), 25|26|28|29|30|31|43 => Pixel_t'(X"6",X"7",X"7"), 32|33|34|35 => Pixel_t'(X"7",X"7",X"7"), 36|37 => Pixel_t'(X"7",X"8",X"8"), 38|39 => Pixel_t'(X"8",X"8",X"8"), 40 => Pixel_t'(X"9",X"9",X"9"), 42 => Pixel_t'(X"a",X"9",X"9"), 41 => Pixel_t'(X"b",X"b",X"b")),
    -- 20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 25 => Pixel_t'(X"1",X"2",X"1"), 45 => Pixel_t'(X"2",X"3",X"3"), 26 => Pixel_t'(X"3",X"3",X"3"), 27|28|44 => Pixel_t'(X"3",X"4",X"4"), 29|43 => Pixel_t'(X"4",X"4",X"4"), 30|31 => Pixel_t'(X"4",X"5",X"5"), 42 => Pixel_t'(X"4",X"5",X"6"), 32|33 => Pixel_t'(X"5",X"5",X"5"), 34|35|36 => Pixel_t'(X"5",X"6",X"6"), 41 => Pixel_t'(X"6",X"6",X"6"), 38 => Pixel_t'(X"6",X"6",X"8"), 37|39 => Pixel_t'(X"6",X"7",X"8"), 40 => Pixel_t'(X"7",X"7",X"7")),
    -- 21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 27|28|45 => Pixel_t'(X"1",X"1",X"1"), 29|30|31 => Pixel_t'(X"2",X"2",X"2"), 32 => Pixel_t'(X"2",X"3",X"3"), 33 => Pixel_t'(X"3",X"3",X"3"), 34 => Pixel_t'(X"3",X"3",X"4"), 35|44 => Pixel_t'(X"3",X"4",X"4"), 36|42 => Pixel_t'(X"4",X"4",X"4"), 43 => Pixel_t'(X"4",X"4",X"5"), 41 => Pixel_t'(X"4",X"5",X"5"), 37|38 => Pixel_t'(X"4",X"5",X"6"), 39 => Pixel_t'(X"5",X"5",X"7"), 40 => Pixel_t'(X"5",X"6",X"6")),
    -- 22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 32|33|34|44 => Pixel_t'(X"1",X"1",X"1"), 35 => Pixel_t'(X"2",X"2",X"2"), 36 => Pixel_t'(X"2",X"3",X"3"), 37|41|42 => Pixel_t'(X"3",X"3",X"3"), 38 => Pixel_t'(X"3",X"4",X"3"), 39|40|43 => Pixel_t'(X"4",X"4",X"4")),
    -- 23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0"), 40 => Pixel_t'(X"1",X"1",X"0"), 39 => Pixel_t'(X"1",X"1",X"1"), 37|38 => Pixel_t'(X"2",X"2",X"2")),
    -- 24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"0",X"0",X"0")));



    -- SCORE --------------------------------------------------------------------------------------------------------------------------

    constant score_9 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|10|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|10|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|13|14 => Pixel_t'("00","00","00"), 9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_8 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_7 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|3|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_6 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 2|3|4|5 => Pixel_t'("11","11","11")),
        2 => (0|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3|4 => Pixel_t'("11","11","11")),
        3 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        11 => (0|4|13|14 => Pixel_t'("00","00","00"), 1|2|3|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|4|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_5 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|11|14 => Pixel_t'("00","00","00"), 1|2|3|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|11|12|14 => Pixel_t'("00","00","00"), 1|2|3|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_4 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 2|3|11|12 => Pixel_t'("11","11","11")),
        2 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_3 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_2 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|11|12|14 => Pixel_t'("00","00","00"), 1|2|3|13 => Pixel_t'("11","11","11")),
        20 => (0|4|5|6|7|8|9|10|11|14 => Pixel_t'("00","00","00"), 1|2|3|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_1 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|2|3|4|5|11|12|13|14 => Pixel_t'("00","00","00"), 6|7|8|9|10 => Pixel_t'("11","11","11")),
        2 => (0|1|2|11|12|13|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10 => Pixel_t'("11","11","11")),
        3 => (0|1|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 2|3|4|8|9|10 => Pixel_t'("11","11","11")),
        4 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        5 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        11 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_0 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|10|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|10|14 => Pixel_t'("00","00","00"), 1|2|3|9|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|4|5|6|7|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|8|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|4|5|6|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|7|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|4|5|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|6|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|5|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|4|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

end package;