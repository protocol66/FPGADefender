library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.my_data_types.all;

package bitmaps is
    constant line_sizeX : positive := 640;
    constant line_sizeY : positive := 2;

    constant ship_sizeX : positive := 25;
    constant ship_sizeY : positive := 25;

    constant score_sizeX : positive := 100;
    constant score_sizeY : positive := 100;


    constant H_LINE : bit_map_t (0 to line_sizeY-1, 0 to line_sizeX-1) := (others => (others => WHITE));
    constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) := (others => (others => TEAL));




    constant score_bit_test : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
   

    (0 => (48|60 => Pixel_t'(X"3",X"4",X"3"), 75 => Pixel_t'(X"4",X"5",X"3"), 26|76 => Pixel_t'(X"4",X"5",X"4"), 27|61 => Pixel_t'(X"4",X"6",X"3"), 49 => Pixel_t'(X"5",X"5",X"5"), 47|62 => Pixel_t'(X"6",X"8",X"5"), 30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|65|67|68|69|70|71 => Pixel_t'(X"6",X"9",X"4"), 29|45|46|63|64|66|72 => Pixel_t'(X"6",X"9",X"5"), 59 => Pixel_t'(X"7",X"7",X"7"), 74 => Pixel_t'(X"7",X"8",X"5"), 28|73 => Pixel_t'(X"7",X"9",X"5"), 25 => Pixel_t'(X"b",X"b",X"c"), 50|77 => Pixel_t'(X"b",X"c",X"c"), 58 => Pixel_t'(X"c",X"c",X"c"), 0|20|21|22|23|52|53|54|55|79|80|81|82|83|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 24|51|56|57|78 => Pixel_t'(X"e",X"e",X"f")),
    1 => (58 => Pixel_t'(X"3",X"4",X"3"), 77 => Pixel_t'(X"3",X"4",X"4"), 25 => Pixel_t'(X"3",X"5",X"3"), 50 => Pixel_t'(X"4",X"4",X"4"), 59 => Pixel_t'(X"4",X"6",X"3"), 49 => Pixel_t'(X"5",X"6",X"4"), 26|76 => Pixel_t'(X"5",X"7",X"4"), 60 => Pixel_t'(X"6",X"8",X"5"), 28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"6",X"9",X"4"), 27|47|61|62|74|75 => Pixel_t'(X"6",X"9",X"5"), 57 => Pixel_t'(X"7",X"8",X"8"), 48 => Pixel_t'(X"7",X"9",X"5"), 51 => Pixel_t'(X"9",X"a",X"a"), 24 => Pixel_t'(X"a",X"a",X"b"), 78 => Pixel_t'(X"b",X"b",X"c"), 56 => Pixel_t'(X"c",X"c",X"d"), 0|16|17|18|19|20|21|22|54|80|81|82|83|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 53 => Pixel_t'(X"e",X"d",X"f"), 23|52|55|79 => Pixel_t'(X"e",X"e",X"f")),
    2 => (24|51 => Pixel_t'(X"3",X"4",X"3"), 78 => Pixel_t'(X"4",X"4",X"4"), 56 => Pixel_t'(X"4",X"5",X"4"), 57 => Pixel_t'(X"4",X"6",X"4"), 77 => Pixel_t'(X"5",X"7",X"5"), 25|50|58 => Pixel_t'(X"6",X"8",X"5"), 27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|61|62|63|64|65|66|67|68|69|70|71|72|73|74 => Pixel_t'(X"6",X"9",X"4"), 60|75|76 => Pixel_t'(X"6",X"9",X"5"), 52 => Pixel_t'(X"7",X"7",X"7"), 26|49|59 => Pixel_t'(X"7",X"9",X"5"), 55 => Pixel_t'(X"9",X"9",X"9"), 23 => Pixel_t'(X"9",X"9",X"a"), 79 => Pixel_t'(X"b",X"c",X"d"), 18|53|54 => Pixel_t'(X"d",X"d",X"e"), 0|16|17|19|20|21|81|82|83|84 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 22|80 => Pixel_t'(X"e",X"e",X"f")),
    3 => (23 => Pixel_t'(X"3",X"4",X"3"), 55 => Pixel_t'(X"3",X"5",X"3"), 52 => Pixel_t'(X"4",X"5",X"3"), 79 => Pixel_t'(X"4",X"5",X"5"), 53|54 => Pixel_t'(X"5",X"6",X"5"), 78 => Pixel_t'(X"5",X"7",X"4"), 24|56 => Pixel_t'(X"6",X"8",X"5"), 26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76 => Pixel_t'(X"6",X"9",X"4"), 50|58 => Pixel_t'(X"6",X"9",X"5"), 25|51|57|77 => Pixel_t'(X"7",X"9",X"5"), 22 => Pixel_t'(X"9",X"a",X"a"), 80 => Pixel_t'(X"d",X"d",X"e"), 0|16|17|19|20|82|83|84 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|18|81|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 21 => Pixel_t'(X"e",X"e",X"f")),
    4 => (22 => Pixel_t'(X"3",X"4",X"3"), 53|54 => Pixel_t'(X"3",X"5",X"3"), 79 => Pixel_t'(X"4",X"6",X"3"), 23 => Pixel_t'(X"6",X"8",X"5"), 25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77 => Pixel_t'(X"6",X"9",X"4"), 49|50|51|56|57|58 => Pixel_t'(X"6",X"9",X"5"), 80 => Pixel_t'(X"7",X"8",X"8"), 24 => Pixel_t'(X"7",X"9",X"4"), 52|78 => Pixel_t'(X"7",X"9",X"5"), 55 => Pixel_t'(X"7",X"9",X"6"), 21 => Pixel_t'(X"a",X"b",X"b"), 0|16|17|18|19|83|84 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|82|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 20|81 => Pixel_t'(X"e",X"e",X"f")),
    5 => (80 => Pixel_t'(X"3",X"4",X"3"), 54 => Pixel_t'(X"3",X"5",X"2"), 21 => Pixel_t'(X"3",X"5",X"3"), 55 => Pixel_t'(X"6",X"8",X"4"), 22|53|79 => Pixel_t'(X"6",X"8",X"5"), 23|24|25|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|47|48|49|50|51|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|77|78 => Pixel_t'(X"6",X"9",X"4"), 26|45|46|52|76 => Pixel_t'(X"6",X"9",X"5"), 20|81 => Pixel_t'(X"b",X"c",X"c"), 0|15|16|17|18|83|84|85 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|82|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 19 => Pixel_t'(X"e",X"e",X"f")),
    6 => (55 => Pixel_t'(X"4",X"6",X"3"), 20 => Pixel_t'(X"4",X"6",X"5"), 80 => Pixel_t'(X"5",X"6",X"4"), 21|54 => Pixel_t'(X"5",X"7",X"4"), 23|24|25|26|27|28|29|30|31|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|77|78 => Pixel_t'(X"6",X"9",X"4"), 22|32|76 => Pixel_t'(X"6",X"9",X"5"), 81 => Pixel_t'(X"7",X"7",X"8"), 53|56|79 => Pixel_t'(X"7",X"9",X"5"), 15|19 => Pixel_t'(X"d",X"d",X"e"), 0|14|16|17|83|84 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 18 => Pixel_t'(X"e",X"d",X"f"), 82 => Pixel_t'(X"e",X"e",X"f")),
    7 => (55 => Pixel_t'(X"3",X"5",X"2"), 81 => Pixel_t'(X"4",X"5",X"4"), 20 => Pixel_t'(X"4",X"6",X"3"), 54|56|80 => Pixel_t'(X"6",X"8",X"5"), 22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|45|46|47|48|49|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'(X"6",X"9",X"4"), 37|38|39|40|41|42|43|44|57 => Pixel_t'(X"6",X"9",X"5"), 19 => Pixel_t'(X"7",X"7",X"7"), 21 => Pixel_t'(X"7",X"9",X"5"), 82 => Pixel_t'(X"c",X"c",X"d"), 0|13|14|15|16|17|84 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|85|86|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 18|83 => Pixel_t'(X"e",X"e",X"f")),
    8 => (40|41|42 => Pixel_t'(X"3",X"5",X"3"), 39 => Pixel_t'(X"3",X"6",X"3"), 19 => Pixel_t'(X"4",X"5",X"3"), 38|43|56 => Pixel_t'(X"4",X"6",X"3"), 44|55|81 => Pixel_t'(X"4",X"6",X"4"), 37|45 => Pixel_t'(X"5",X"7",X"4"), 36|46 => Pixel_t'(X"6",X"8",X"5"), 21|22|23|24|25|26|27|28|29|30|31|32|33|50|51|52|53|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'(X"6",X"9",X"4"), 20|34|35|47|49 => Pixel_t'(X"6",X"9",X"5"), 48|54|57|80 => Pixel_t'(X"7",X"9",X"5"), 82 => Pixel_t'(X"9",X"9",X"9"), 18 => Pixel_t'(X"a",X"b",X"b"), 0|14|15|16|84|85|86 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|87|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 17|83 => Pixel_t'(X"e",X"e",X"f")),
    9 => (35|36|46|47|56 => Pixel_t'(X"3",X"5",X"2"), 45 => Pixel_t'(X"3",X"5",X"3"), 18 => Pixel_t'(X"4",X"5",X"4"), 37|44 => Pixel_t'(X"4",X"6",X"3"), 38|48 => Pixel_t'(X"4",X"6",X"4"), 34 => Pixel_t'(X"4",X"7",X"4"), 82 => Pixel_t'(X"5",X"6",X"6"), 39|40|41|42|43 => Pixel_t'(X"5",X"7",X"4"), 81 => Pixel_t'(X"6",X"7",X"4"), 19|33|49|55 => Pixel_t'(X"6",X"8",X"5"), 21|22|23|24|25|26|27|28|29|30|52|53|54|58|59|60|61|62|63|64|65|66|67|68|69|70|72|73|74|75|77|78|79|80 => Pixel_t'(X"6",X"9",X"4"), 20|31|32|50|51|57|71|76 => Pixel_t'(X"6",X"9",X"5"), 17 => Pixel_t'(X"c",X"d",X"e"), 0|15|84|85|86|87 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|16|83|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f")),
    10 => (33|49 => Pixel_t'(X"3",X"5",X"2"), 50|56 => Pixel_t'(X"3",X"5",X"3"), 82 => Pixel_t'(X"4",X"5",X"4"), 18|32|34|48 => Pixel_t'(X"4",X"6",X"3"), 35|47|51|57 => Pixel_t'(X"5",X"8",X"4"), 31 => Pixel_t'(X"6",X"8",X"5"), 20|21|23|24|25|26|27|28|39|40|54|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80 => Pixel_t'(X"6",X"9",X"4"), 22|29|30|36|37|41|42|43|44|45|46|53|55 => Pixel_t'(X"6",X"9",X"5"), 17 => Pixel_t'(X"7",X"8",X"8"), 19|38|52|81 => Pixel_t'(X"7",X"9",X"5"), 83 => Pixel_t'(X"c",X"c",X"d"), 0|13|14|15|85|86|87 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|88|89|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 16|84 => Pixel_t'(X"e",X"e",X"f")),
    11 => (31 => Pixel_t'(X"2",X"5",X"2"), 51 => Pixel_t'(X"3",X"5",X"2"), 17|52 => Pixel_t'(X"3",X"5",X"3"), 32 => Pixel_t'(X"4",X"6",X"3"), 30|82 => Pixel_t'(X"4",X"6",X"4"), 50|56|57 => Pixel_t'(X"4",X"7",X"4"), 18|33|49|53 => Pixel_t'(X"6",X"8",X"5"), 19|20|21|27|28|36|37|38|39|40|41|42|43|44|45|46|59|60|61|76|77|78|79|80 => Pixel_t'(X"6",X"9",X"4"), 22|23|24|25|26|29|34|35|47|54|62|63|64|65|66|67|68|69|70|71|72|73|74|75 => Pixel_t'(X"6",X"9",X"5"), 48|55|58|81 => Pixel_t'(X"7",X"9",X"5"), 83 => Pixel_t'(X"a",X"a",X"b"), 16 => Pixel_t'(X"c",X"c",X"d"), 0|13|85|86|87|88|89 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 14 => Pixel_t'(X"e",X"d",X"f"), 15|84 => Pixel_t'(X"e",X"e",X"f")),
    12 => (53 => Pixel_t'(X"2",X"5",X"2"), 29|71|72|73|74 => Pixel_t'(X"3",X"5",X"2"), 30|66|67|68|69|70|75 => Pixel_t'(X"3",X"5",X"3"), 65 => Pixel_t'(X"3",X"6",X"3"), 57|64|76 => Pixel_t'(X"4",X"6",X"3"), 54 => Pixel_t'(X"4",X"6",X"4"), 52 => Pixel_t'(X"4",X"7",X"3"), 63 => Pixel_t'(X"4",X"7",X"4"), 17 => Pixel_t'(X"5",X"6",X"4"), 82 => Pixel_t'(X"5",X"7",X"5"), 62 => Pixel_t'(X"5",X"8",X"4"), 16 => Pixel_t'(X"6",X"7",X"7"), 56|79 => Pixel_t'(X"6",X"8",X"4"), 28|31|61|77 => Pixel_t'(X"6",X"8",X"5"), 19|20|21|26|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49 => Pixel_t'(X"6",X"9",X"4"), 18|22|23|24|25|33|50|51|59|60|78|80 => Pixel_t'(X"6",X"9",X"5"), 27|32|55|81 => Pixel_t'(X"7",X"9",X"5"), 58 => Pixel_t'(X"7",X"9",X"6"), 83 => Pixel_t'(X"8",X"9",X"9"), 0|13|14|85|86|87|88|89 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|9|10|11|12|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 15|84 => Pixel_t'(X"e",X"e",X"f")),
    13 => (57 => Pixel_t'(X"3",X"4",X"2"), 28|60|61|62|77|78|79|80 => Pixel_t'(X"3",X"5",X"2"), 55 => Pixel_t'(X"3",X"5",X"3"), 54|59 => Pixel_t'(X"3",X"6",X"3"), 16 => Pixel_t'(X"4",X"5",X"3"), 83 => Pixel_t'(X"4",X"5",X"5"), 63|76 => Pixel_t'(X"4",X"6",X"3"), 58|64|82 => Pixel_t'(X"4",X"6",X"4"), 27|29|65|66|75|81 => Pixel_t'(X"5",X"7",X"4"), 56 => Pixel_t'(X"6",X"7",X"5"), 67 => Pixel_t'(X"6",X"8",X"4"), 53|68|69|70|71|72|73|74 => Pixel_t'(X"6",X"8",X"5"), 18|19|20|21|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51 => Pixel_t'(X"6",X"9",X"4"), 17|22|23|24|25|26|31 => Pixel_t'(X"6",X"9",X"5"), 30|52 => Pixel_t'(X"7",X"9",X"5"), 15 => Pixel_t'(X"b",X"c",X"c"), 84 => Pixel_t'(X"c",X"c",X"c"), 0|8|9|13|87|88|89 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|10|11|12|90|91|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 14|85|86 => Pixel_t'(X"e",X"e",X"f")),
    14 => (56|57 => Pixel_t'(X"2",X"3",X"2"), 84 => Pixel_t'(X"3",X"4",X"3"), 82 => Pixel_t'(X"3",X"5",X"3"), 27 => Pixel_t'(X"3",X"6",X"2"), 83 => Pixel_t'(X"4",X"5",X"3"), 81 => Pixel_t'(X"4",X"6",X"3"), 58 => Pixel_t'(X"4",X"6",X"4"), 16 => Pixel_t'(X"5",X"6",X"4"), 85 => Pixel_t'(X"5",X"6",X"6"), 55|59 => Pixel_t'(X"5",X"7",X"4"), 80 => Pixel_t'(X"5",X"8",X"4"), 15 => Pixel_t'(X"6",X"7",X"7"), 26|28|60 => Pixel_t'(X"6",X"8",X"4"), 78 => Pixel_t'(X"6",X"8",X"5"), 18|19|20|21|22|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|52|65|66|67|68|69|70|71|72|73|74|75 => Pixel_t'(X"6",X"9",X"4"), 17|23|24|25|50|51|53|61|62|63|64|76|77|79 => Pixel_t'(X"6",X"9",X"5"), 54 => Pixel_t'(X"7",X"9",X"5"), 86 => Pixel_t'(X"a",X"a",X"a"), 87 => Pixel_t'(X"d",X"d",X"e"), 0|8|9|10|13|89|91 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|11|12|90|92|93|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 14|88 => Pixel_t'(X"e",X"e",X"f")),
    15 => (57 => Pixel_t'(X"3",X"5",X"3"), 15|86 => Pixel_t'(X"4",X"5",X"3"), 87 => Pixel_t'(X"4",X"5",X"4"), 85 => Pixel_t'(X"5",X"7",X"4"), 56|84 => Pixel_t'(X"6",X"8",X"5"), 58 => Pixel_t'(X"6",X"8",X"6"), 17|19|20|21|22|23|24|25|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|53|54|60|63|64|65|66|67|68|69|70|71|72|73|77|78|79|80 => Pixel_t'(X"6",X"9",X"4"), 16|18|26|27|50|51|52|61|62|74|75|76|81|82 => Pixel_t'(X"6",X"9",X"5"), 55|59|83 => Pixel_t'(X"7",X"9",X"5"), 88 => Pixel_t'(X"9",X"a",X"a"), 14 => Pixel_t'(X"c",X"c",X"d"), 0|9|10|11|91|92|93 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|12|13|89|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 90 => Pixel_t'(X"e",X"e",X"f")),
    16 => (58 => Pixel_t'(X"3",X"5",X"2"), 88 => Pixel_t'(X"3",X"5",X"3"), 15 => Pixel_t'(X"4",X"6",X"3"), 89 => Pixel_t'(X"5",X"6",X"6"), 57 => Pixel_t'(X"5",X"7",X"4"), 87 => Pixel_t'(X"5",X"7",X"5"), 59 => Pixel_t'(X"6",X"8",X"4"), 17|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|42|43|44|45|46|47|48|49|50|51|52|53|54|55|61|62|63|64|65|66|67|68|73|74|77|78|79|80|81|82|83|84 => Pixel_t'(X"6",X"9",X"4"), 16|18|41|56|60|69|70|71|72|75|76|85 => Pixel_t'(X"6",X"9",X"5"), 14 => Pixel_t'(X"7",X"8",X"8"), 86 => Pixel_t'(X"7",X"9",X"5"), 90 => Pixel_t'(X"c",X"d",X"d"), 0|9|10|11|92|93 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|7|8|12|94|95|96|97|98|99 => Pixel_t'(X"d",X"e",X"f"), 13|91 => Pixel_t'(X"e",X"e",X"f")),
    17 => (59 => Pixel_t'(X"3",X"5",X"2"), 90 => Pixel_t'(X"4",X"5",X"4"), 14 => Pixel_t'(X"4",X"5",X"5"), 89 => Pixel_t'(X"4",X"6",X"4"), 58 => Pixel_t'(X"5",X"7",X"5"), 15|60 => Pixel_t'(X"6",X"8",X"5"), 16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|42|43|44|52|62|63|64|65|66|67|68|72|73|74|75|76|81|82|83|84|85|86 => Pixel_t'(X"6",X"9",X"4"), 41|45|46|47|48|49|50|51|53|54|55|56|69|70|71|77|78|79|80|87|88 => Pixel_t'(X"6",X"9",X"5"), 61 => Pixel_t'(X"7",X"9",X"5"), 57 => Pixel_t'(X"7",X"9",X"6"), 91 => Pixel_t'(X"b",X"b",X"c"), 11|13 => Pixel_t'(X"d",X"d",X"e"), 0|4|5|6|7|8|9|10|93|94|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|12|95|96 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    18 => (60 => Pixel_t'(X"2",X"4",X"2"), 48|49|50|51|52|53|54|55 => Pixel_t'(X"3",X"5",X"2"), 56 => Pixel_t'(X"3",X"5",X"3"), 47 => Pixel_t'(X"3",X"6",X"3"), 91 => Pixel_t'(X"4",X"4",X"4"), 14 => Pixel_t'(X"4",X"5",X"3"), 59 => Pixel_t'(X"4",X"5",X"4"), 57 => Pixel_t'(X"4",X"6",X"3"), 46 => Pixel_t'(X"4",X"6",X"4"), 58 => Pixel_t'(X"5",X"6",X"5"), 45 => Pixel_t'(X"5",X"7",X"4"), 90 => Pixel_t'(X"5",X"7",X"5"), 80 => Pixel_t'(X"5",X"8",X"4"), 79|81 => Pixel_t'(X"6",X"8",X"4"), 44|61|78|82|83 => Pixel_t'(X"6",X"8",X"5"), 16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|63|64|65|66|67|68|71 => Pixel_t'(X"6",X"9",X"4"), 41|43|62|69|70|72|73|77|84|86|87|88 => Pixel_t'(X"6",X"9",X"5"), 15|42|74|75|76|85|89 => Pixel_t'(X"7",X"9",X"5"), 13 => Pixel_t'(X"a",X"a",X"b"), 92 => Pixel_t'(X"b",X"b",X"c"), 0|4|5|6|7|8|9|10|11|94|97|98 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|95|96|99 => Pixel_t'(X"d",X"e",X"f"), 12|93 => Pixel_t'(X"e",X"e",X"f")),
    19 => (60 => Pixel_t'(X"1",X"3",X"1"), 61 => Pixel_t'(X"2",X"4",X"1"), 44|78|79|80 => Pixel_t'(X"2",X"5",X"2"), 92 => Pixel_t'(X"3",X"4",X"4"), 43|45|76|77|81|82|83|84|85 => Pixel_t'(X"3",X"5",X"2"), 59|86 => Pixel_t'(X"3",X"5",X"3"), 75 => Pixel_t'(X"3",X"6",X"3"), 42|46|58|74|87 => Pixel_t'(X"4",X"6",X"3"), 14|47|56|57|73|88 => Pixel_t'(X"5",X"7",X"4"), 62 => Pixel_t'(X"5",X"7",X"5"), 13 => Pixel_t'(X"6",X"6",X"6"), 91 => Pixel_t'(X"6",X"7",X"6"), 48|55|89 => Pixel_t'(X"6",X"8",X"4"), 41|49|50|51|52|53|54 => Pixel_t'(X"6",X"8",X"5"), 16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|64|65|66|67|68 => Pixel_t'(X"6",X"9",X"4"), 39|63|69|70|71|72 => Pixel_t'(X"6",X"9",X"5"), 15 => Pixel_t'(X"7",X"9",X"4"), 40|90 => Pixel_t'(X"7",X"9",X"5"), 93 => Pixel_t'(X"b",X"b",X"c"), 0|4|5|6|7|8|9|10|95|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|11|96 => Pixel_t'(X"d",X"e",X"f"), 12|94 => Pixel_t'(X"e",X"e",X"f")),
    20 => (90 => Pixel_t'(X"3",X"4",X"2"), 92 => Pixel_t'(X"3",X"4",X"3"), 41|62|72|73|89 => Pixel_t'(X"3",X"5",X"2"), 40|71|88 => Pixel_t'(X"3",X"5",X"3"), 13 => Pixel_t'(X"4",X"5",X"4"), 42|74|87 => Pixel_t'(X"4",X"6",X"3"), 91 => Pixel_t'(X"4",X"6",X"4"), 39|61|63|70|75|86 => Pixel_t'(X"5",X"7",X"4"), 43 => Pixel_t'(X"5",X"8",X"4"), 49|50|51|69|76|85 => Pixel_t'(X"6",X"8",X"4"), 14|48|52|53|84 => Pixel_t'(X"6",X"8",X"5"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|36|65 => Pixel_t'(X"6",X"9",X"4"), 35|37|38|44|54|60|64|66|67|77|78|82|83 => Pixel_t'(X"6",X"9",X"5"), 45|47|55|56|57|58|59|68|79|81 => Pixel_t'(X"7",X"9",X"5"), 46|80 => Pixel_t'(X"7",X"9",X"6"), 93 => Pixel_t'(X"9",X"9",X"a"), 12 => Pixel_t'(X"c",X"c",X"d"), 0|7|8|9|10|96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|6|95 => Pixel_t'(X"d",X"e",X"f"), 11|94 => Pixel_t'(X"e",X"e",X"f")),
    21 => (53 => Pixel_t'(X"2",X"4",X"2"), 48|52|54 => Pixel_t'(X"3",X"4",X"2"), 93 => Pixel_t'(X"3",X"4",X"3"), 38|39|47|49|50|51|55|69 => Pixel_t'(X"3",X"5",X"2"), 63|68 => Pixel_t'(X"3",X"5",X"3"), 46|92 => Pixel_t'(X"4",X"5",X"3"), 13|56|70|81|82 => Pixel_t'(X"4",X"6",X"3"), 64|79|80 => Pixel_t'(X"4",X"6",X"4"), 40|45|57|67|71|78|83|84|85|91 => Pixel_t'(X"5",X"7",X"4"), 77 => Pixel_t'(X"5",X"7",X"5"), 37 => Pixel_t'(X"6",X"8",X"4"), 44|58|62|72|76|86|87|90 => Pixel_t'(X"6",X"8",X"5"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35 => Pixel_t'(X"6",X"9",X"4"), 14|41|59|60|66 => Pixel_t'(X"6",X"9",X"5"), 94 => Pixel_t'(X"7",X"8",X"8"), 36|42|61|65|73|74|75|88|89 => Pixel_t'(X"7",X"9",X"5"), 43 => Pixel_t'(X"7",X"9",X"6"), 12 => Pixel_t'(X"a",X"a",X"b"), 95 => Pixel_t'(X"d",X"d",X"e"), 0|6|7|8|9|10|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|5|96 => Pixel_t'(X"d",X"e",X"f"), 11 => Pixel_t'(X"e",X"e",X"f")),
    22 => (37|44|58|59|66|74|75|76|77|85|86|87|88 => Pixel_t'(X"3",X"5",X"2"), 43|64|67 => Pixel_t'(X"3",X"5",X"3"), 45 => Pixel_t'(X"3",X"6",X"3"), 94 => Pixel_t'(X"4",X"5",X"4"), 56|57|60|73|78|79|80|81|82|83|84|89 => Pixel_t'(X"4",X"6",X"3"), 65 => Pixel_t'(X"4",X"6",X"4"), 95 => Pixel_t'(X"5",X"6",X"5"), 13|36|38|42|46|55|68|72|90 => Pixel_t'(X"5",X"7",X"4"), 12 => Pixel_t'(X"6",X"7",X"7"), 47|61 => Pixel_t'(X"6",X"8",X"4"), 48|53|54|71 => Pixel_t'(X"6",X"8",X"5"), 15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'(X"6",X"9",X"4"), 14|34|39|41|49|50|51|52 => Pixel_t'(X"6",X"9",X"5"), 91 => Pixel_t'(X"7",X"8",X"5"), 63|93 => Pixel_t'(X"7",X"8",X"6"), 35|40|62 => Pixel_t'(X"7",X"9",X"5"), 69|70|92 => Pixel_t'(X"7",X"9",X"6"), 6|96 => Pixel_t'(X"d",X"d",X"e"), 0|5|7|8|98|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|4|11|97 => Pixel_t'(X"d",X"e",X"f"), 9|10 => Pixel_t'(X"e",X"e",X"f")),
    23 => (12 => Pixel_t'(X"2",X"3",X"2"), 64 => Pixel_t'(X"2",X"4",X"2"), 36|41|42|61|62|70|71|72|91 => Pixel_t'(X"3",X"5",X"2"), 65|90 => Pixel_t'(X"3",X"5",X"3"), 95 => Pixel_t'(X"4",X"5",X"4"), 35|51|52|60|69|73|89|92 => Pixel_t'(X"4",X"6",X"3"), 50 => Pixel_t'(X"4",X"7",X"3"), 11 => Pixel_t'(X"5",X"5",X"5"), 53 => Pixel_t'(X"5",X"7",X"3"), 43|47|48|49|74 => Pixel_t'(X"5",X"7",X"4"), 63 => Pixel_t'(X"5",X"7",X"5"), 54|80|88 => Pixel_t'(X"5",X"8",X"4"), 40 => Pixel_t'(X"6",X"7",X"4"), 81|82|83 => Pixel_t'(X"6",X"8",X"4"), 13|34|37|55|59|66|68|75|79|87|93 => Pixel_t'(X"6",X"8",X"5"), 14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|84 => Pixel_t'(X"6",X"9",X"4"), 33|44|45|46|56|76|78|85|86 => Pixel_t'(X"6",X"9",X"5"), 96 => Pixel_t'(X"7",X"7",X"7"), 38|39|57|77 => Pixel_t'(X"7",X"9",X"5"), 58|67|94 => Pixel_t'(X"7",X"9",X"6"), 10 => Pixel_t'(X"8",X"8",X"8"), 9 => Pixel_t'(X"c",X"d",X"d"), 0|4|5|6|7|98 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|99 => Pixel_t'(X"d",X"e",X"f"), 8|97 => Pixel_t'(X"e",X"e",X"f")),
    24 => (63 => Pixel_t'(X"3",X"4",X"2"), 34|40|67|68|93 => Pixel_t'(X"3",X"5",X"2"), 12|94 => Pixel_t'(X"3",X"5",X"3"), 10 => Pixel_t'(X"4",X"5",X"3"), 9 => Pixel_t'(X"4",X"5",X"4"), 35|39|57|64|66|69|86 => Pixel_t'(X"4",X"6",X"3"), 82 => Pixel_t'(X"4",X"6",X"4"), 92 => Pixel_t'(X"4",X"7",X"4"), 96 => Pixel_t'(X"5",X"5",X"5"), 44|81|83|85 => Pixel_t'(X"5",X"6",X"4"), 88 => Pixel_t'(X"5",X"7",X"3"), 33|41|56|70|77|87 => Pixel_t'(X"5",X"7",X"4"), 11|45|62|78 => Pixel_t'(X"5",X"7",X"5"), 58|76 => Pixel_t'(X"5",X"8",X"4"), 43 => Pixel_t'(X"6",X"7",X"4"), 79|80|84|95 => Pixel_t'(X"6",X"7",X"5"), 46 => Pixel_t'(X"6",X"7",X"6"), 38|42|59|65|71|89|91 => Pixel_t'(X"6",X"8",X"5"), 14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'(X"6",X"9",X"4"), 13|30|31|32|36|75 => Pixel_t'(X"6",X"9",X"5"), 37|60|61|72|73|74|90 => Pixel_t'(X"7",X"9",X"5"), 55 => Pixel_t'(X"8",X"9",X"7"), 47|54 => Pixel_t'(X"8",X"9",X"8"), 53 => Pixel_t'(X"9",X"a",X"9"), 8 => Pixel_t'(X"9",X"a",X"a"), 52 => Pixel_t'(X"b",X"b",X"a"), 48 => Pixel_t'(X"c",X"c",X"c"), 49|51 => Pixel_t'(X"c",X"d",X"c"), 50 => Pixel_t'(X"d",X"d",X"d"), 97 => Pixel_t'(X"d",X"d",X"e"), 0|4|5|6|99 => Pixel_t'(X"d",X"d",X"f"), 1|2|3|98 => Pixel_t'(X"d",X"e",X"f"), 7 => Pixel_t'(X"e",X"e",X"f")),
    25 => (82 => Pixel_t'(X"1",X"0",X"1"), 80|81|83 => Pixel_t'(X"1",X"1",X"1"), 79 => Pixel_t'(X"2",X"2",X"2"), 95 => Pixel_t'(X"2",X"4",X"2"), 8 => Pixel_t'(X"3",X"4",X"3"), 32|33|38 => Pixel_t'(X"3",X"5",X"2"), 48 => Pixel_t'(X"4",X"3",X"4"), 47|49|96 => Pixel_t'(X"4",X"4",X"4"), 60 => Pixel_t'(X"4",X"5",X"3"), 12|31|39|42|65|66|74|90 => Pixel_t'(X"4",X"6",X"3"), 46|78|84 => Pixel_t'(X"5",X"5",X"5"), 59|75 => Pixel_t'(X"5",X"6",X"4"), 37|41|61|94 => Pixel_t'(X"5",X"7",X"4"), 30|67|91 => Pixel_t'(X"5",X"8",X"4"), 50 => Pixel_t'(X"6",X"6",X"6"), 89 => Pixel_t'(X"6",X"7",X"5"), 76 => Pixel_t'(X"6",X"7",X"6"), 9|73 => Pixel_t'(X"6",X"8",X"4"), 11|34|40|62 => Pixel_t'(X"6",X"8",X"5"), 14|15|16|17|18|19|20|21|22|23|24|25|26|70|71 => Pixel_t'(X"6",X"9",X"4"), 13|27|28|29|68|69|72|93 => Pixel_t'(X"6",X"9",X"5"), 58 => Pixel_t'(X"7",X"7",X"6"), 77 => Pixel_t'(X"7",X"7",X"7"), 64 => Pixel_t'(X"7",X"8",X"5"), 88 => Pixel_t'(X"7",X"8",X"7"), 10|35|36|63|92 => Pixel_t'(X"7",X"9",X"5"), 7|45 => Pixel_t'(X"8",X"8",X"8"), 43 => Pixel_t'(X"9",X"a",X"9"), 57 => Pixel_t'(X"a",X"a",X"9"), 87 => Pixel_t'(X"a",X"b",X"a"), 44|85 => Pixel_t'(X"b",X"b",X"b"), 51 => Pixel_t'(X"b",X"b",X"c"), 86 => Pixel_t'(X"d",X"d",X"d"), 97 => Pixel_t'(X"d",X"d",X"e"), 0|2|3|4|5|99 => Pixel_t'(X"d",X"d",X"f"), 1 => Pixel_t'(X"d",X"e",X"f"), 56 => Pixel_t'(X"e",X"e",X"e"), 6|98 => Pixel_t'(X"e",X"e",X"f"), 52|53|54|55 => Pixel_t'(X"f",X"f",X"f")),
    26 => (47|48|49|50|51|80|81|82|83|84 => Pixel_t'(X"0",X"0",X"0"), 77 => Pixel_t'(X"1",X"1",X"1"), 46 => Pixel_t'(X"1",X"1",X"2"), 44|45|85 => Pixel_t'(X"2",X"2",X"2"), 29 => Pixel_t'(X"2",X"5",X"2"), 78 => Pixel_t'(X"3",X"3",X"3"), 92 => Pixel_t'(X"3",X"4",X"2"), 96 => Pixel_t'(X"3",X"4",X"3"), 30|37 => Pixel_t'(X"3",X"5",X"2"), 7 => Pixel_t'(X"3",X"5",X"3"), 62|63 => Pixel_t'(X"4",X"5",X"3"), 12|31|36|72 => Pixel_t'(X"4",X"6",X"3"), 28 => Pixel_t'(X"4",X"7",X"3"), 40 => Pixel_t'(X"5",X"6",X"5"), 97 => Pixel_t'(X"5",X"6",X"6"), 11|64 => Pixel_t'(X"5",X"7",X"4"), 79 => Pixel_t'(X"6",X"6",X"6"), 38|39 => Pixel_t'(X"6",X"7",X"5"), 73|91 => Pixel_t'(X"6",X"7",X"6"), 71 => Pixel_t'(X"6",X"8",X"4"), 32|35|93|95 => Pixel_t'(X"6",X"8",X"5"), 9|14|15|16|17|18|19|20|21|22|23|24|25|26|67|68|69 => Pixel_t'(X"6",X"9",X"4"), 8|10|13|27|65|70|94 => Pixel_t'(X"6",X"9",X"5"), 52 => Pixel_t'(X"7",X"7",X"7"), 61 => Pixel_t'(X"7",X"8",X"7"), 33|34|66 => Pixel_t'(X"7",X"9",X"5"), 76 => Pixel_t'(X"8",X"8",X"9"), 6 => Pixel_t'(X"8",X"9",X"9"), 41 => Pixel_t'(X"9",X"9",X"8"), 43|74 => Pixel_t'(X"a",X"b",X"a"), 60 => Pixel_t'(X"b",X"c",X"b"), 86 => Pixel_t'(X"c",X"c",X"d"), 90 => Pixel_t'(X"c",X"d",X"c"), 98 => Pixel_t'(X"d",X"d",X"e"), 0|2|3|4 => Pixel_t'(X"d",X"d",X"f"), 42 => Pixel_t'(X"d",X"e",X"d"), 1 => Pixel_t'(X"d",X"e",X"f"), 75 => Pixel_t'(X"e",X"e",X"e"), 5|99 => Pixel_t'(X"e",X"e",X"f"), 59 => Pixel_t'(X"e",X"f",X"e"), 89 => Pixel_t'(X"f",X"f",X"e"), 53|54|55|56|57|58|87|88 => Pixel_t'(X"f",X"f",X"f")),
    27 => (43|44|47|48|49|50|51|52|76|77|81|82|83|84|85 => Pixel_t'(X"0",X"0",X"0"), 80 => Pixel_t'(X"2",X"2",X"2"), 35 => Pixel_t'(X"2",X"5",X"2"), 86 => Pixel_t'(X"3",X"3",X"3"), 6|93 => Pixel_t'(X"3",X"4",X"3"), 65 => Pixel_t'(X"3",X"5",X"2"), 94 => Pixel_t'(X"4",X"5",X"3"), 34 => Pixel_t'(X"4",X"6",X"3"), 11|36|97 => Pixel_t'(X"4",X"6",X"4"), 70 => Pixel_t'(X"5",X"6",X"3"), 38 => Pixel_t'(X"5",X"6",X"4"), 12|95 => Pixel_t'(X"5",X"7",X"4"), 64 => Pixel_t'(X"6",X"6",X"5"), 98 => Pixel_t'(X"6",X"6",X"7"), 37 => Pixel_t'(X"6",X"7",X"5"), 28|29 => Pixel_t'(X"6",X"8",X"4"), 7|33 => Pixel_t'(X"6",X"8",X"5"), 9|14|15|16|17|18|19|20|21|22|23|24|25|26|27|67|68 => Pixel_t'(X"6",X"9",X"4"), 8|10|13|66|69 => Pixel_t'(X"6",X"9",X"5"), 92 => Pixel_t'(X"7",X"7",X"6"), 71|96 => Pixel_t'(X"7",X"8",X"6"), 30|31|32 => Pixel_t'(X"7",X"9",X"5"), 53 => Pixel_t'(X"8",X"8",X"8"), 39 => Pixel_t'(X"9",X"a",X"9"), 75 => Pixel_t'(X"a",X"a",X"a"), 42 => Pixel_t'(X"b",X"a",X"a"), 5|63|72|78 => Pixel_t'(X"b",X"b",X"b"), 45|46 => Pixel_t'(X"c",X"c",X"c"), 99 => Pixel_t'(X"d",X"d",X"e"), 0|2|3 => Pixel_t'(X"d",X"d",X"f"), 1 => Pixel_t'(X"d",X"e",X"f"), 40 => Pixel_t'(X"e",X"e",X"e"), 4 => Pixel_t'(X"e",X"e",X"f"), 62 => Pixel_t'(X"f",X"f",X"e"), 41|54|55|56|57|58|59|60|61|73|74|79|87|88|89|90|91 => Pixel_t'(X"f",X"f",X"f")),
    28 => (43|44|47|48|51|52|76|77|80|81|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 49 => Pixel_t'(X"1",X"0",X"1"), 50|53 => Pixel_t'(X"1",X"1",X"1"), 42|82 => Pixel_t'(X"2",X"2",X"2"), 75 => Pixel_t'(X"3",X"3",X"3"), 33 => Pixel_t'(X"3",X"5",X"2"), 78 => Pixel_t'(X"4",X"3",X"4"), 83 => Pixel_t'(X"4",X"4",X"4"), 98 => Pixel_t'(X"4",X"4",X"5"), 32|96 => Pixel_t'(X"4",X"5",X"3"), 11|34|66 => Pixel_t'(X"4",X"6",X"3"), 5 => Pixel_t'(X"5",X"6",X"5"), 6|31|36|69 => Pixel_t'(X"5",X"7",X"4"), 97 => Pixel_t'(X"5",X"7",X"5"), 12 => Pixel_t'(X"5",X"8",X"4"), 37 => Pixel_t'(X"6",X"7",X"5"), 29|30|35|68 => Pixel_t'(X"6",X"8",X"5"), 8|9|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 10|24|25|26|27|28 => Pixel_t'(X"6",X"9",X"5"), 79 => Pixel_t'(X"7",X"7",X"7"), 95 => Pixel_t'(X"7",X"8",X"7"), 7|67 => Pixel_t'(X"7",X"9",X"5"), 45 => Pixel_t'(X"8",X"8",X"9"), 65 => Pixel_t'(X"9",X"9",X"8"), 46 => Pixel_t'(X"9",X"9",X"9"), 70 => Pixel_t'(X"a",X"a",X"9"), 87 => Pixel_t'(X"a",X"a",X"a"), 94 => Pixel_t'(X"b",X"b",X"b"), 99 => Pixel_t'(X"c",X"c",X"d"), 38 => Pixel_t'(X"c",X"d",X"c"), 4|54 => Pixel_t'(X"d",X"d",X"e"), 0|2|3 => Pixel_t'(X"d",X"d",X"f"), 1 => Pixel_t'(X"d",X"e",X"f"), 41|93 => Pixel_t'(X"e",X"e",X"e"), 39|40|55|56|57|58|59|60|61|62|63|64|71|72|73|74|88|89|90|91|92 => Pixel_t'(X"f",X"f",X"f")),
    29 => (42|43|44|45|46|47|52|53|75|76|77|78|79|80|85|86 => Pixel_t'(X"0",X"0",X"0"), 81 => Pixel_t'(X"1",X"1",X"1"), 48 => Pixel_t'(X"2",X"2",X"2"), 51 => Pixel_t'(X"3",X"3",X"3"), 26|27|28|29|30 => Pixel_t'(X"3",X"5",X"2"), 11|31 => Pixel_t'(X"3",X"5",X"3"), 87|97 => Pixel_t'(X"4",X"4",X"4"), 5 => Pixel_t'(X"4",X"5",X"3"), 25 => Pixel_t'(X"4",X"7",X"3"), 66 => Pixel_t'(X"5",X"6",X"5"), 32|35 => Pixel_t'(X"5",X"7",X"4"), 98 => Pixel_t'(X"6",X"6",X"6"), 67|68 => Pixel_t'(X"6",X"7",X"5"), 12 => Pixel_t'(X"6",X"8",X"4"), 33 => Pixel_t'(X"6",X"8",X"5"), 7|8|9|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 10|24 => Pixel_t'(X"6",X"9",X"5"), 84 => Pixel_t'(X"7",X"7",X"7"), 6|34 => Pixel_t'(X"7",X"9",X"5"), 54 => Pixel_t'(X"8",X"8",X"8"), 36 => Pixel_t'(X"8",X"9",X"7"), 4 => Pixel_t'(X"9",X"a",X"a"), 41 => Pixel_t'(X"b",X"b",X"b"), 49|74 => Pixel_t'(X"c",X"c",X"c"), 69|96 => Pixel_t'(X"c",X"d",X"c"), 50|82 => Pixel_t'(X"d",X"d",X"d"), 99 => Pixel_t'(X"d",X"d",X"e"), 0|2 => Pixel_t'(X"d",X"d",X"f"), 1 => Pixel_t'(X"d",X"e",X"f"), 3 => Pixel_t'(X"e",X"e",X"f"), 37 => Pixel_t'(X"f",X"f",X"e"), 38|39|40|55|56|57|58|59|60|61|62|63|64|65|70|71|72|73|83|88|89|90|91|92|93|94|95 => Pixel_t'(X"f",X"f",X"f")),
    30 => (42|43|44|45|46|47|52|53|75|76|77|78|80|85|86 => Pixel_t'(X"0",X"0",X"0"), 79|81 => Pixel_t'(X"0",X"0",X"1"), 87 => Pixel_t'(X"2",X"1",X"2"), 48 => Pixel_t'(X"3",X"3",X"3"), 25 => Pixel_t'(X"3",X"5",X"2"), 11 => Pixel_t'(X"3",X"5",X"3"), 67 => Pixel_t'(X"4",X"4",X"3"), 54 => Pixel_t'(X"4",X"4",X"4"), 4 => Pixel_t'(X"4",X"5",X"4"), 51|98 => Pixel_t'(X"5",X"5",X"5"), 34 => Pixel_t'(X"5",X"7",X"4"), 84 => Pixel_t'(X"6",X"6",X"6"), 5|27|28 => Pixel_t'(X"6",X"8",X"4"), 12|24|26 => Pixel_t'(X"6",X"8",X"5"), 6|7|8|9|13|14|15|16|17|18|19|20|21|22 => Pixel_t'(X"6",X"9",X"4"), 10|23|29|30|33 => Pixel_t'(X"6",X"9",X"5"), 66 => Pixel_t'(X"7",X"7",X"7"), 31|32 => Pixel_t'(X"7",X"9",X"5"), 41 => Pixel_t'(X"8",X"8",X"8"), 74 => Pixel_t'(X"a",X"a",X"a"), 35 => Pixel_t'(X"b",X"b",X"a"), 97 => Pixel_t'(X"b",X"b",X"b"), 82 => Pixel_t'(X"c",X"c",X"c"), 68 => Pixel_t'(X"d",X"d",X"d"), 3|99 => Pixel_t'(X"d",X"d",X"e"), 0 => Pixel_t'(X"d",X"d",X"f"), 1|2 => Pixel_t'(X"d",X"e",X"f"), 88 => Pixel_t'(X"e",X"e",X"e"), 36|37|38|39|40|49|50|55|56|57|58|59|60|61|62|63|64|65|69|70|71|72|73|83|89|90|91|92|93|94|95|96 => Pixel_t'(X"f",X"f",X"f")),
    31 => (42|43|44|47|48|51|52|53|75|76|77|81|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 80|87 => Pixel_t'(X"1",X"1",X"1"), 82 => Pixel_t'(X"2",X"2",X"2"), 54 => Pixel_t'(X"3",X"3",X"3"), 78 => Pixel_t'(X"3",X"3",X"4"), 25 => Pixel_t'(X"3",X"5",X"2"), 11 => Pixel_t'(X"3",X"5",X"3"), 45 => Pixel_t'(X"4",X"4",X"4"), 4 => Pixel_t'(X"4",X"5",X"3"), 33 => Pixel_t'(X"4",X"6",X"4"), 83 => Pixel_t'(X"5",X"4",X"5"), 98 => Pixel_t'(X"5",X"5",X"6"), 10|24|26 => Pixel_t'(X"6",X"8",X"5"), 6|7|8|9|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 12|28|30|31|32 => Pixel_t'(X"6",X"9",X"5"), 41|49|66 => Pixel_t'(X"7",X"7",X"7"), 46|50 => Pixel_t'(X"7",X"7",X"8"), 5|27|29 => Pixel_t'(X"7",X"9",X"5"), 74 => Pixel_t'(X"9",X"9",X"9"), 3 => Pixel_t'(X"9",X"9",X"a"), 34 => Pixel_t'(X"a",X"b",X"a"), 79|99 => Pixel_t'(X"b",X"b",X"c"), 67 => Pixel_t'(X"c",X"c",X"c"), 88 => Pixel_t'(X"d",X"d",X"d"), 1 => Pixel_t'(X"d",X"d",X"e"), 0 => Pixel_t'(X"d",X"d",X"f"), 2 => Pixel_t'(X"e",X"e",X"f"), 35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|65|68|69|70|71|72|73|89|90|91|92|93|94|95|96|97 => Pixel_t'(X"f",X"f",X"f")),
    32 => (42|43|44|47|48|49|50|51|52|53|75|76|77|80|81|82|83|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 87 => Pixel_t'(X"0",X"0",X"1"), 78 => Pixel_t'(X"2",X"1",X"2"), 54 => Pixel_t'(X"2",X"2",X"2"), 26 => Pixel_t'(X"3",X"5",X"2"), 27 => Pixel_t'(X"3",X"5",X"3"), 11|28 => Pixel_t'(X"3",X"6",X"3"), 29 => Pixel_t'(X"4",X"6",X"3"), 3 => Pixel_t'(X"4",X"6",X"4"), 25 => Pixel_t'(X"4",X"7",X"4"), 45|79 => Pixel_t'(X"5",X"5",X"5"), 32 => Pixel_t'(X"5",X"6",X"4"), 30|31 => Pixel_t'(X"5",X"7",X"4"), 41 => Pixel_t'(X"6",X"6",X"6"), 10 => Pixel_t'(X"6",X"8",X"4"), 4 => Pixel_t'(X"6",X"8",X"5"), 5|6|7|8|9|13|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 12|14|24 => Pixel_t'(X"6",X"9",X"5"), 46|66|74|98 => Pixel_t'(X"8",X"8",X"8"), 99 => Pixel_t'(X"a",X"9",X"a"), 33 => Pixel_t'(X"b",X"b",X"a"), 1|2 => Pixel_t'(X"c",X"d",X"e"), 88 => Pixel_t'(X"d",X"c",X"d"), 0 => Pixel_t'(X"d",X"e",X"f"), 55|65 => Pixel_t'(X"e",X"e",X"e"), 34|35|36|37|38|39|40|56|57|58|59|60|61|62|63|64|67|68|69|70|71|72|73|89|90|91|92|93|94|95|96|97 => Pixel_t'(X"f",X"f",X"f")),
    33 => (42|43|44|45|46|47|48|49|50|51|52|53|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 87 => Pixel_t'(X"1",X"1",X"1"), 31 => Pixel_t'(X"2",X"3",X"1"), 54 => Pixel_t'(X"3",X"3",X"3"), 41 => Pixel_t'(X"4",X"4",X"4"), 3 => Pixel_t'(X"4",X"5",X"3"), 30 => Pixel_t'(X"4",X"6",X"3"), 29 => Pixel_t'(X"5",X"6",X"4"), 32 => Pixel_t'(X"5",X"6",X"5"), 27|28 => Pixel_t'(X"5",X"7",X"4"), 98 => Pixel_t'(X"6",X"6",X"7"), 11 => Pixel_t'(X"6",X"8",X"4"), 26 => Pixel_t'(X"6",X"8",X"5"), 5|6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'(X"6",X"9",X"4"), 25 => Pixel_t'(X"6",X"9",X"5"), 74 => Pixel_t'(X"7",X"7",X"7"), 4 => Pixel_t'(X"7",X"9",X"5"), 2 => Pixel_t'(X"9",X"9",X"a"), 66 => Pixel_t'(X"a",X"a",X"a"), 99 => Pixel_t'(X"a",X"a",X"b"), 65 => Pixel_t'(X"c",X"c",X"c"), 1 => Pixel_t'(X"d",X"d",X"e"), 0 => Pixel_t'(X"d",X"d",X"f"), 88 => Pixel_t'(X"e",X"e",X"e"), 33|34|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|67|68|69|70|71|72|73|89|90|91|92|93|94|95|96|97 => Pixel_t'(X"f",X"f",X"f")),
    34 => (42|43|44|45|46|47|48|49|50|51|52|53|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 87 => Pixel_t'(X"2",X"2",X"2"), 54 => Pixel_t'(X"4",X"4",X"4"), 98 => Pixel_t'(X"4",X"4",X"5"), 32 => Pixel_t'(X"4",X"5",X"3"), 2|41 => Pixel_t'(X"5",X"5",X"5"), 3 => Pixel_t'(X"5",X"7",X"4"), 31 => Pixel_t'(X"6",X"8",X"5"), 4|5|6|7|8|9|10|12|13|14|15|16|17|18|19|20|21|22|23|24|25 => Pixel_t'(X"6",X"9",X"4"), 11|26|27|28|29|30 => Pixel_t'(X"6",X"9",X"5"), 74 => Pixel_t'(X"8",X"8",X"8"), 33 => Pixel_t'(X"9",X"9",X"9"), 65|97 => Pixel_t'(X"a",X"a",X"a"), 66 => Pixel_t'(X"c",X"c",X"c"), 99 => Pixel_t'(X"c",X"c",X"d"), 1 => Pixel_t'(X"c",X"d",X"e"), 0 => Pixel_t'(X"d",X"e",X"f"), 88 => Pixel_t'(X"f",X"e",X"e"), 34|35|36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|67|68|69|70|71|72|73|89|90|91|92|93|94|95|96 => Pixel_t'(X"f",X"f",X"f")),
    35 => (42|43|44|45|46|47|48|49|50|51|52|53|75|76|77|78|79|80|81|82|83|84|85|86 => Pixel_t'(X"0",X"0",X"0"), 97 => Pixel_t'(X"3",X"3",X"4"), 2 => Pixel_t'(X"3",X"5",X"3"), 33 => Pixel_t'(X"4",X"5",X"3"), 32 => Pixel_t'(X"6",X"8",X"5"), 4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'(X"6",X"9",X"4"), 3|31 => Pixel_t'(X"6",X"9",X"5"), 34|65 => Pixel_t'(X"7",X"8",X"7"), 41|87 => Pixel_t'(X"8",X"8",X"8"), 54 => Pixel_t'(X"9",X"9",X"9"), 96 => Pixel_t'(X"a",X"a",X"a"), 1|74 => Pixel_t'(X"b",X"b",X"b"), 98 => Pixel_t'(X"b",X"b",X"c"), 99 => Pixel_t'(X"d",X"d",X"e"), 35|66 => Pixel_t'(X"e",X"e",X"e"), 0 => Pixel_t'(X"e",X"e",X"f"), 36|37|38|39|40|55|56|57|58|59|60|61|62|63|64|67|68|69|70|71|72|73|88|89|90|91|92|93|94|95 => Pixel_t'(X"f",X"f",X"f")),
    36 => (42|43|44|45|46|47|48|49|50|51|52|76|77|78|79|80|81|82|83|84|85 => Pixel_t'(X"0",X"0",X"0"), 96 => Pixel_t'(X"3",X"3",X"3"), 53|65|75 => Pixel_t'(X"4",X"4",X"4"), 35 => Pixel_t'(X"4",X"5",X"4"), 95 => Pixel_t'(X"5",X"5",X"4"), 86 => Pixel_t'(X"5",X"5",X"5"), 2 => Pixel_t'(X"5",X"7",X"4"), 34 => Pixel_t'(X"5",X"7",X"5"), 64 => Pixel_t'(X"6",X"6",X"6"), 4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32 => Pixel_t'(X"6",X"9",X"4"), 3|33 => Pixel_t'(X"6",X"9",X"5"), 1 => Pixel_t'(X"7",X"7",X"7"), 94 => Pixel_t'(X"9",X"9",X"9"), 36 => Pixel_t'(X"a",X"a",X"a"), 97 => Pixel_t'(X"b",X"b",X"c"), 41 => Pixel_t'(X"c",X"c",X"c"), 63|93 => Pixel_t'(X"d",X"d",X"d"), 98 => Pixel_t'(X"d",X"d",X"e"), 99 => Pixel_t'(X"d",X"e",X"f"), 0 => Pixel_t'(X"e",X"e",X"f"), 54 => Pixel_t'(X"f",X"e",X"f"), 37|38|39|40|55|56|57|58|59|60|61|62|66|67|68|69|70|71|72|73|74|87|88|89|90|91|92 => Pixel_t'(X"f",X"f",X"f")),
    37 => (43|44|45|46|47|48|49|50|51|77|78|79|80|81|82|83|84 => Pixel_t'(X"0",X"0",X"0"), 76 => Pixel_t'(X"2",X"1",X"2"), 52 => Pixel_t'(X"3",X"3",X"3"), 63 => Pixel_t'(X"3",X"4",X"3"), 93 => Pixel_t'(X"3",X"5",X"3"), 65 => Pixel_t'(X"4",X"4",X"3"), 85 => Pixel_t'(X"4",X"4",X"4"), 36|94 => Pixel_t'(X"4",X"5",X"3"), 1 => Pixel_t'(X"4",X"5",X"4"), 92|96 => Pixel_t'(X"5",X"5",X"5"), 64 => Pixel_t'(X"5",X"6",X"5"), 37 => Pixel_t'(X"6",X"6",X"5"), 66 => Pixel_t'(X"6",X"6",X"6"), 95 => Pixel_t'(X"6",X"7",X"5"), 2|35 => Pixel_t'(X"6",X"8",X"5"), 3|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'(X"6",X"9",X"4"), 4 => Pixel_t'(X"6",X"9",X"5"), 62 => Pixel_t'(X"7",X"8",X"7"), 34 => Pixel_t'(X"7",X"9",X"5"), 42|91 => Pixel_t'(X"8",X"8",X"8"), 97 => Pixel_t'(X"b",X"b",X"c"), 38 => Pixel_t'(X"b",X"c",X"b"), 90 => Pixel_t'(X"c",X"c",X"c"), 0 => Pixel_t'(X"c",X"c",X"d"), 67 => Pixel_t'(X"c",X"d",X"c"), 75 => Pixel_t'(X"d",X"d",X"d"), 98 => Pixel_t'(X"d",X"d",X"e"), 99 => Pixel_t'(X"d",X"e",X"f"), 61 => Pixel_t'(X"e",X"e",X"d"), 53|89 => Pixel_t'(X"e",X"e",X"e"), 39|40|41|54|55|56|57|58|59|60|68|69|70|71|72|73|74|86|87|88 => Pixel_t'(X"f",X"f",X"f")),
    38 => (45|46|47|48|49|79|80|82 => Pixel_t'(X"0",X"0",X"0"), 81 => Pixel_t'(X"0",X"0",X"1"), 44|50|83 => Pixel_t'(X"1",X"1",X"1"), 78 => Pixel_t'(X"2",X"2",X"2"), 66 => Pixel_t'(X"2",X"4",X"2"), 90 => Pixel_t'(X"3",X"4",X"3"), 38|67 => Pixel_t'(X"4",X"5",X"3"), 96 => Pixel_t'(X"4",X"5",X"5"), 1|91 => Pixel_t'(X"4",X"6",X"3"), 65 => Pixel_t'(X"4",X"6",X"4"), 68|89 => Pixel_t'(X"5",X"5",X"4"), 51|77|84 => Pixel_t'(X"5",X"5",X"5"), 62|95 => Pixel_t'(X"5",X"6",X"4"), 39|61|88 => Pixel_t'(X"5",X"6",X"5"), 32 => Pixel_t'(X"5",X"7",X"3"), 33 => Pixel_t'(X"5",X"7",X"4"), 69|87 => Pixel_t'(X"6",X"6",X"6"), 92 => Pixel_t'(X"6",X"7",X"4"), 37 => Pixel_t'(X"6",X"7",X"5"), 3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'(X"6",X"9",X"4"), 31 => Pixel_t'(X"6",X"9",X"5"), 43 => Pixel_t'(X"7",X"7",X"7"), 63 => Pixel_t'(X"7",X"8",X"5"), 60|86 => Pixel_t'(X"7",X"8",X"7"), 2 => Pixel_t'(X"7",X"9",X"4"), 34|35|36|93 => Pixel_t'(X"7",X"9",X"5"), 64|94 => Pixel_t'(X"7",X"9",X"6"), 70 => Pixel_t'(X"8",X"8",X"7"), 85 => Pixel_t'(X"8",X"9",X"8"), 0 => Pixel_t'(X"8",X"9",X"9"), 40|59|71 => Pixel_t'(X"a",X"a",X"a"), 72 => Pixel_t'(X"c",X"c",X"c"), 76|97 => Pixel_t'(X"c",X"c",X"d"), 98 => Pixel_t'(X"c",X"d",X"e"), 52 => Pixel_t'(X"d",X"d",X"d"), 99 => Pixel_t'(X"d",X"e",X"f"), 73 => Pixel_t'(X"e",X"e",X"d"), 58 => Pixel_t'(X"e",X"e",X"e"), 74 => Pixel_t'(X"f",X"e",X"f"), 41|42|53|54|55|56|57|75 => Pixel_t'(X"f",X"f",X"f")),
    39 => (82 => Pixel_t'(X"2",X"3",X"2"), 79 => Pixel_t'(X"3",X"3",X"3"), 81|83|94 => Pixel_t'(X"3",X"4",X"3"), 33|65 => Pixel_t'(X"3",X"5",X"2"), 34 => Pixel_t'(X"3",X"6",X"3"), 58|80 => Pixel_t'(X"4",X"4",X"3"), 40|59|72|84|85 => Pixel_t'(X"4",X"5",X"3"), 0|73 => Pixel_t'(X"4",X"5",X"4"), 71|86 => Pixel_t'(X"4",X"6",X"3"), 41 => Pixel_t'(X"5",X"5",X"4"), 57|74 => Pixel_t'(X"5",X"5",X"5"), 70 => Pixel_t'(X"5",X"6",X"3"), 95 => Pixel_t'(X"5",X"6",X"6"), 60|69|87|93 => Pixel_t'(X"5",X"7",X"4"), 32 => Pixel_t'(X"5",X"8",X"4"), 75|78 => Pixel_t'(X"6",X"6",X"5"), 46 => Pixel_t'(X"6",X"6",X"7"), 39 => Pixel_t'(X"6",X"7",X"4"), 1|35 => Pixel_t'(X"6",X"8",X"4"), 61|64|66|68|88|89 => Pixel_t'(X"6",X"8",X"5"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'(X"6",X"9",X"4"), 31|36|63|91 => Pixel_t'(X"6",X"9",X"5"), 47 => Pixel_t'(X"7",X"7",X"7"), 37|38|62|67|90|92 => Pixel_t'(X"7",X"9",X"5"), 48|76 => Pixel_t'(X"8",X"8",X"8"), 56 => Pixel_t'(X"8",X"9",X"8"), 45 => Pixel_t'(X"9",X"8",X"9"), 42|77 => Pixel_t'(X"9",X"9",X"8"), 49 => Pixel_t'(X"9",X"9",X"9"), 44|55 => Pixel_t'(X"c",X"c",X"c"), 96 => Pixel_t'(X"c",X"c",X"d"), 98 => Pixel_t'(X"c",X"c",X"e"), 50 => Pixel_t'(X"d",X"c",X"d"), 43 => Pixel_t'(X"d",X"d",X"d"), 97 => Pixel_t'(X"d",X"d",X"e"), 99 => Pixel_t'(X"e",X"d",X"f"), 54 => Pixel_t'(X"e",X"e",X"e"), 53 => Pixel_t'(X"e",X"e",X"f"), 51|52 => Pixel_t'(X"f",X"f",X"f")),
    40 => (35|64 => Pixel_t'(X"3",X"5",X"2"), 0 => Pixel_t'(X"3",X"5",X"3"), 36 => Pixel_t'(X"3",X"6",X"3"), 43|44|54|55 => Pixel_t'(X"4",X"5",X"3"), 45|50 => Pixel_t'(X"4",X"5",X"4"), 42|56 => Pixel_t'(X"4",X"6",X"3"), 92 => Pixel_t'(X"4",X"6",X"4"), 34 => Pixel_t'(X"4",X"7",X"4"), 46|51 => Pixel_t'(X"5",X"5",X"4"), 48|49 => Pixel_t'(X"5",X"5",X"5"), 53 => Pixel_t'(X"5",X"6",X"4"), 47|52|93 => Pixel_t'(X"5",X"6",X"5"), 57|65|79 => Pixel_t'(X"5",X"7",X"4"), 37|76 => Pixel_t'(X"5",X"8",X"4"), 78 => Pixel_t'(X"6",X"7",X"4"), 75|77|80|81 => Pixel_t'(X"6",X"8",X"4"), 41|58|63|74|82 => Pixel_t'(X"6",X"8",X"5"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|67|89|90 => Pixel_t'(X"6",X"9",X"4"), 1|32|33|38|61|62|66|68|69|70|71|72|73|84|85|86|87|88|91 => Pixel_t'(X"6",X"9",X"5"), 39|40|59|60|83 => Pixel_t'(X"7",X"9",X"5"), 94 => Pixel_t'(X"a",X"a",X"b"), 97|98 => Pixel_t'(X"d",X"d",X"e"), 99 => Pixel_t'(X"d",X"d",X"f"), 95 => Pixel_t'(X"d",X"e",X"f"), 96 => Pixel_t'(X"e",X"e",X"f")),
    41 => (37|38|63 => Pixel_t'(X"3",X"5",X"2"), 92 => Pixel_t'(X"4",X"5",X"4"), 39 => Pixel_t'(X"4",X"7",X"3"), 36 => Pixel_t'(X"4",X"7",X"4"), 0|47|48|49|50|51|62|64 => Pixel_t'(X"5",X"7",X"4"), 40|44|45|46|52|53|60|61|91 => Pixel_t'(X"6",X"8",X"5"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|57|66|67|68|69|70|73|74|75|76|77|81|82|83|84|85|86|87|88|89|90 => Pixel_t'(X"6",X"9",X"4"), 1|33|34|35|54|55|56|58|59|65|71|72|78|79|80 => Pixel_t'(X"6",X"9",X"5"), 41|42|43 => Pixel_t'(X"7",X"9",X"5"), 93 => Pixel_t'(X"d",X"d",X"e"), 96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 95 => Pixel_t'(X"e",X"d",X"f"), 94 => Pixel_t'(X"e",X"e",X"f")),
    42 => (40|60|61|62 => Pixel_t'(X"3",X"5",X"2"), 39|41 => Pixel_t'(X"3",X"5",X"3"), 59 => Pixel_t'(X"3",X"6",X"3"), 42 => Pixel_t'(X"4",X"6",X"3"), 91 => Pixel_t'(X"4",X"6",X"4"), 38|58 => Pixel_t'(X"5",X"7",X"4"), 43 => Pixel_t'(X"5",X"8",X"4"), 63 => Pixel_t'(X"6",X"8",X"4"), 44|57 => Pixel_t'(X"6",X"8",X"5"), 2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 1|37|45|46|47|48|49|50|51|52|53|54|55|56|65|90 => Pixel_t'(X"6",X"9",X"5"), 92 => Pixel_t'(X"7",X"8",X"8"), 0|36|64 => Pixel_t'(X"7",X"9",X"5"), 94|95|96|97|99 => Pixel_t'(X"d",X"d",X"f"), 98 => Pixel_t'(X"d",X"e",X"f"), 93 => Pixel_t'(X"e",X"e",X"f")),
    43 => (43|44|45|46|47|48|49|50|51|57 => Pixel_t'(X"3",X"5",X"2"), 52|53|54|55|56|58 => Pixel_t'(X"3",X"5",X"3"), 42 => Pixel_t'(X"4",X"6",X"3"), 91 => Pixel_t'(X"5",X"5",X"5"), 41|59|90 => Pixel_t'(X"5",X"7",X"4"), 40|60 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88 => Pixel_t'(X"6",X"9",X"4"), 38|39|61|62 => Pixel_t'(X"6",X"9",X"5"), 0 => Pixel_t'(X"7",X"9",X"4"), 89 => Pixel_t'(X"7",X"9",X"5"), 92 => Pixel_t'(X"d",X"d",X"e"), 93|94|95|96|99 => Pixel_t'(X"d",X"d",X"f"), 97|98 => Pixel_t'(X"d",X"e",X"f")),
    44 => (90 => Pixel_t'(X"4",X"5",X"5"), 89 => Pixel_t'(X"4",X"6",X"4"), 53|54|55 => Pixel_t'(X"5",X"8",X"4"), 48|49|50|56 => Pixel_t'(X"6",X"8",X"4"), 45|46|47|51|52|57|58 => Pixel_t'(X"6",X"8",X"5"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|37|38|39|40|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|81|83|84|85|86 => Pixel_t'(X"6",X"9",X"4"), 36|41|42|43|44|59|60|79|80|82|87 => Pixel_t'(X"6",X"9",X"5"), 88 => Pixel_t'(X"7",X"9",X"5"), 91 => Pixel_t'(X"c",X"c",X"d"), 93|94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    45 => (58 => Pixel_t'(X"3",X"5",X"2"), 88 => Pixel_t'(X"4",X"5",X"3"), 57 => Pixel_t'(X"4",X"6",X"3"), 89 => Pixel_t'(X"5",X"6",X"6"), 56|59|86|87 => Pixel_t'(X"6",X"8",X"5"), 0|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|53|61|62|63|64|65|66|67|70|71|72|73|74|77|78|79|80|81 => Pixel_t'(X"6",X"9",X"4"), 1|45|46|47|48|49|50|51|52|60|68|69|75|76|82|83|84 => Pixel_t'(X"6",X"9",X"5"), 54|55|85 => Pixel_t'(X"7",X"9",X"5"), 90 => Pixel_t'(X"c",X"c",X"d"), 92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 91 => Pixel_t'(X"e",X"e",X"f")),
    46 => (55 => Pixel_t'(X"3",X"5",X"3"), 86 => Pixel_t'(X"4",X"5",X"4"), 56|68|69 => Pixel_t'(X"4",X"6",X"3"), 85 => Pixel_t'(X"4",X"6",X"4"), 57 => Pixel_t'(X"5",X"7",X"4"), 54|58 => Pixel_t'(X"6",X"8",X"4"), 70|84 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|48|49|50|51|59|60|61|62|63|64|65|66|67|73|74|75|76|78|79|80 => Pixel_t'(X"6",X"9",X"4"), 0|7|44|45|46|47|52|72|77|81|82|83 => Pixel_t'(X"6",X"9",X"5"), 53|71 => Pixel_t'(X"7",X"9",X"5"), 87 => Pixel_t'(X"8",X"9",X"9"), 88 => Pixel_t'(X"b",X"b",X"c"), 89 => Pixel_t'(X"d",X"d",X"e"), 91|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 90|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    47 => (85 => Pixel_t'(X"2",X"3",X"2"), 84 => Pixel_t'(X"2",X"4",X"2"), 70 => Pixel_t'(X"3",X"4",X"2"), 54|83 => Pixel_t'(X"3",X"5",X"2"), 53|69|71|82 => Pixel_t'(X"4",X"6",X"3"), 55 => Pixel_t'(X"5",X"7",X"3"), 81 => Pixel_t'(X"5",X"7",X"4"), 52 => Pixel_t'(X"5",X"8",X"4"), 72|80 => Pixel_t'(X"6",X"8",X"4"), 68|79 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|46|47|48|58|59|60|61|62|63|64|65|66|67 => Pixel_t'(X"6",X"9",X"4"), 0|5|6|44|45|49|50|51|56|73|75|76|77|78 => Pixel_t'(X"6",X"9",X"5"), 57|74 => Pixel_t'(X"7",X"9",X"5"), 86 => Pixel_t'(X"b",X"b",X"b"), 89|90|91|99 => Pixel_t'(X"d",X"d",X"f"), 92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 87|88 => Pixel_t'(X"e",X"e",X"f")),
    48 => (73 => Pixel_t'(X"2",X"4",X"2"), 78 => Pixel_t'(X"2",X"5",X"2"), 74 => Pixel_t'(X"3",X"4",X"2"), 51|52|72|75|76|77|79|80 => Pixel_t'(X"3",X"5",X"2"), 71|81 => Pixel_t'(X"4",X"6",X"3"), 85 => Pixel_t'(X"4",X"6",X"4"), 82 => Pixel_t'(X"4",X"7",X"3"), 53 => Pixel_t'(X"4",X"7",X"4"), 50 => Pixel_t'(X"5",X"7",X"4"), 83 => Pixel_t'(X"5",X"8",X"4"), 86 => Pixel_t'(X"6",X"6",X"6"), 70 => Pixel_t'(X"6",X"8",X"4"), 84 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|46|47|55|56|57|61|62|63|64|65|66|67 => Pixel_t'(X"6",X"9",X"4"), 0|5|6|44|45|48|49|54|58|59|60|68 => Pixel_t'(X"6",X"9",X"5"), 69 => Pixel_t'(X"7",X"9",X"5"), 87 => Pixel_t'(X"d",X"d",X"e"), 89|90|99 => Pixel_t'(X"d",X"d",X"f"), 91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 88 => Pixel_t'(X"e",X"e",X"f")),
    49 => (74 => Pixel_t'(X"2",X"3",X"1"), 49|50 => Pixel_t'(X"3",X"5",X"2"), 86 => Pixel_t'(X"4",X"5",X"3"), 75 => Pixel_t'(X"4",X"6",X"3"), 73 => Pixel_t'(X"4",X"6",X"4"), 48|51 => Pixel_t'(X"5",X"7",X"4"), 76|77 => Pixel_t'(X"5",X"8",X"4"), 87 => Pixel_t'(X"6",X"7",X"6"), 78 => Pixel_t'(X"6",X"8",X"4"), 47 => Pixel_t'(X"6",X"8",X"5"), 1|3|4|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|79|83|84 => Pixel_t'(X"6",X"9",X"4"), 0|2|5|6|44|45|46|52|53|54|72|80|81|82|85 => Pixel_t'(X"6",X"9",X"5"), 88 => Pixel_t'(X"d",X"d",X"e"), 89|90|99 => Pixel_t'(X"d",X"d",X"f"), 91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    50 => (47 => Pixel_t'(X"3",X"5",X"2"), 75 => Pixel_t'(X"3",X"6",X"2"), 46 => Pixel_t'(X"3",X"6",X"3"), 87 => Pixel_t'(X"4",X"5",X"3"), 48 => Pixel_t'(X"4",X"6",X"3"), 49 => Pixel_t'(X"5",X"7",X"4"), 45|74|76 => Pixel_t'(X"6",X"8",X"4"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|77|78|79|80|81|82|83|84|85 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|44|50|51|72|73|86 => Pixel_t'(X"6",X"9",X"5"), 88 => Pixel_t'(X"7",X"8",X"8"), 90|91|99 => Pixel_t'(X"d",X"d",X"f"), 89|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    51 => (88 => Pixel_t'(X"3",X"5",X"3"), 46 => Pixel_t'(X"4",X"6",X"3"), 45 => Pixel_t'(X"5",X"8",X"4"), 47 => Pixel_t'(X"6",X"8",X"4"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|72|73|74|75|76|77|78|80|81|82|83|84|85|86 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|44|48|70|71|79|87 => Pixel_t'(X"6",X"9",X"5"), 89 => Pixel_t'(X"9",X"a",X"a"), 91|92|99 => Pixel_t'(X"d",X"d",X"f"), 93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 90 => Pixel_t'(X"e",X"e",X"f")),
    52 => (89 => Pixel_t'(X"4",X"5",X"4"), 88 => Pixel_t'(X"6",X"8",X"5"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|85|86 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|82|83|84|87 => Pixel_t'(X"6",X"9",X"5"), 90 => Pixel_t'(X"c",X"c",X"d"), 92|93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 91 => Pixel_t'(X"e",X"e",X"f")),
    53 => (89 => Pixel_t'(X"4",X"6",X"4"), 90 => Pixel_t'(X"6",X"7",X"7"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|85|86|87 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|82|83|84|88 => Pixel_t'(X"6",X"9",X"5"), 92|93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 91 => Pixel_t'(X"e",X"e",X"f")),
    54 => (90 => Pixel_t'(X"3",X"5",X"3"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|85|86|87|88 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|82|83|84|89 => Pixel_t'(X"6",X"9",X"5"), 91 => Pixel_t'(X"b",X"b",X"c"), 93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    55 => (90 => Pixel_t'(X"5",X"7",X"4"), 1|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|85|86|87|88 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|83|84|89 => Pixel_t'(X"6",X"9",X"5"), 91 => Pixel_t'(X"7",X"7",X"7"), 93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    56 => (91 => Pixel_t'(X"4",X"5",X"4"), 90 => Pixel_t'(X"6",X"8",X"5"), 1|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|32|33|34|35|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|27|28|29|30|31|36|37|38|39 => Pixel_t'(X"6",X"9",X"5"), 92 => Pixel_t'(X"d",X"d",X"e"), 93|94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    57 => (91 => Pixel_t'(X"4",X"5",X"3"), 1|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|32|33|34|35|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|26|27|28|29|30|31|36|37|38|39|90 => Pixel_t'(X"6",X"9",X"5"), 92 => Pixel_t'(X"a",X"a",X"b"), 94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 93 => Pixel_t'(X"e",X"e",X"f")),
    58 => (91 => Pixel_t'(X"5",X"7",X"4"), 1|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|32|33|34|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|26|27|28|29|30|31|35|36|37|38|39|90 => Pixel_t'(X"6",X"9",X"5"), 92 => Pixel_t'(X"7",X"7",X"8"), 94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 93 => Pixel_t'(X"e",X"e",X"f")),
    59 => (92 => Pixel_t'(X"5",X"6",X"5"), 91 => Pixel_t'(X"6",X"8",X"4"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|37|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 0|35|36|38|39|90 => Pixel_t'(X"6",X"9",X"5"), 93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    60 => (92 => Pixel_t'(X"5",X"5",X"5"), 91 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|25|26|27|28|29|30|31|32|37|38|39|40|41|42|43|44|45|46|47|48|49|52|53|54|55|56|58|59|60|64|65|66|67|68|69|70|71|72|73|74|75|76|82|83|84|88|89|90 => Pixel_t'(X"6",X"9",X"4"), 0|23|24|33|34|35|36|50|51|57|61|62|63|77|78|79|80|81|85|86|87 => Pixel_t'(X"6",X"9",X"5"), 93 => Pixel_t'(X"d",X"d",X"e"), 99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    61 => (92 => Pixel_t'(X"4",X"5",X"4"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|25|26|27|28|42|43|44|45|46|47|48|49|52|53|54|55|59|60|64|65|66|67|68|69|70|71|72|73|74|75|76|82|83|84|85|88|89|90 => Pixel_t'(X"6",X"9",X"4"), 0|23|24|29|33|34|35|36|39|40|41|50|51|56|57|58|61|62|63|77|78|79|80|81|86|87|91 => Pixel_t'(X"6",X"9",X"5"), 30|31|32|37|38 => Pixel_t'(X"7",X"9",X"5"), 93 => Pixel_t'(X"c",X"c",X"d"), 99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 94 => Pixel_t'(X"e",X"e",X"f")),
    62 => (34|35 => Pixel_t'(X"4",X"3",X"2"), 36 => Pixel_t'(X"4",X"4",X"2"), 92 => Pixel_t'(X"4",X"4",X"3"), 33 => Pixel_t'(X"5",X"3",X"2"), 37 => Pixel_t'(X"5",X"4",X"2"), 32 => Pixel_t'(X"5",X"4",X"3"), 31|38 => Pixel_t'(X"5",X"5",X"3"), 39 => Pixel_t'(X"5",X"6",X"4"), 30 => Pixel_t'(X"6",X"6",X"4"), 40 => Pixel_t'(X"6",X"7",X"4"), 41|42 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|26|27|46|47|48|49|52|53|54|55|56|58|59|60|64|65|66|67|68|69|70|71|72|73|74|75|76|83|84|85|86|87|88|89 => Pixel_t'(X"6",X"9",X"4"), 0|23|24|25|43|45|50|51|57|61|62|63|77|78|79|80|81|82|90 => Pixel_t'(X"6",X"9",X"5"), 29 => Pixel_t'(X"7",X"8",X"5"), 28|44 => Pixel_t'(X"7",X"9",X"5"), 91 => Pixel_t'(X"7",X"9",X"6"), 93 => Pixel_t'(X"9",X"8",X"8"), 94 => Pixel_t'(X"d",X"d",X"e"), 96|97|99 => Pixel_t'(X"d",X"d",X"f"), 95|98 => Pixel_t'(X"d",X"e",X"f")),
    63 => (42 => Pixel_t'(X"4",X"4",X"2"), 43 => Pixel_t'(X"4",X"5",X"3"), 41|92|93 => Pixel_t'(X"5",X"3",X"2"), 29|91 => Pixel_t'(X"5",X"4",X"2"), 44 => Pixel_t'(X"5",X"6",X"4"), 30|40 => Pixel_t'(X"6",X"3",X"2"), 28|90 => Pixel_t'(X"6",X"7",X"4"), 45 => Pixel_t'(X"6",X"7",X"5"), 46 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|52|53|54|55|56|57|58|59|60|65|66|67|68|69|70|71|72|73|74|75|76|83|84|85|86 => Pixel_t'(X"6",X"9",X"4"), 0|26|27|48|49|50|51|61|62|63|64|77|78|79|80|81|82|87|88 => Pixel_t'(X"6",X"9",X"5"), 39 => Pixel_t'(X"7",X"4",X"2"), 38 => Pixel_t'(X"7",X"4",X"3"), 47|89 => Pixel_t'(X"7",X"9",X"5"), 31 => Pixel_t'(X"8",X"4",X"3"), 37 => Pixel_t'(X"8",X"5",X"3"), 94 => Pixel_t'(X"8",X"7",X"8"), 32 => Pixel_t'(X"9",X"5",X"3"), 33|36 => Pixel_t'(X"9",X"5",X"4"), 34|35 => Pixel_t'(X"9",X"6",X"4"), 96|97|99 => Pixel_t'(X"d",X"d",X"f"), 95|98 => Pixel_t'(X"d",X"e",X"f")),
    64 => (28|45|46 => Pixel_t'(X"5",X"3",X"2"), 47|89 => Pixel_t'(X"5",X"4",X"2"), 94 => Pixel_t'(X"5",X"4",X"3"), 48 => Pixel_t'(X"5",X"5",X"3"), 49|88 => Pixel_t'(X"5",X"6",X"4"), 90 => Pixel_t'(X"6",X"3",X"2"), 27 => Pixel_t'(X"6",X"6",X"4"), 50 => Pixel_t'(X"6",X"7",X"5"), 51|87 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|57|58|59|60|61|66|67|68|69|70|71|72|73|74|75|76|77|81|82|83 => Pixel_t'(X"6",X"9",X"4"), 0|5|6|26|52|53|54|55|56|62|63|64|65|78|79|80|84|85|86 => Pixel_t'(X"6",X"9",X"5"), 44 => Pixel_t'(X"7",X"4",X"2"), 43 => Pixel_t'(X"8",X"5",X"3"), 91 => Pixel_t'(X"9",X"5",X"3"), 29|42 => Pixel_t'(X"9",X"5",X"4"), 30|31|32|33|35|36|37|38|40|41|92 => Pixel_t'(X"a",X"6",X"4"), 93 => Pixel_t'(X"a",X"6",X"5"), 34|39 => Pixel_t'(X"b",X"6",X"4"), 95 => Pixel_t'(X"c",X"c",X"d"), 97|99 => Pixel_t'(X"d",X"d",X"f"), 96|98 => Pixel_t'(X"d",X"e",X"f")),
    65 => (27|50|51|87 => Pixel_t'(X"5",X"3",X"2"), 52 => Pixel_t'(X"5",X"4",X"3"), 53|86 => Pixel_t'(X"5",X"5",X"3"), 54 => Pixel_t'(X"5",X"6",X"4"), 49|88 => Pixel_t'(X"6",X"3",X"2"), 94 => Pixel_t'(X"6",X"4",X"3"), 85 => Pixel_t'(X"6",X"6",X"4"), 26|55 => Pixel_t'(X"6",X"7",X"5"), 56 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79 => Pixel_t'(X"6",X"9",X"4"), 0|6|25|60|61|62|63|64|80|81|82 => Pixel_t'(X"6",X"9",X"5"), 48 => Pixel_t'(X"7",X"4",X"3"), 84 => Pixel_t'(X"7",X"8",X"5"), 57|58|59|83 => Pixel_t'(X"7",X"9",X"5"), 47|89 => Pixel_t'(X"9",X"5",X"3"), 28 => Pixel_t'(X"9",X"6",X"4"), 29|30|31|32|33|34|35|36|37|38|39|40|41|42|44|45|46|90|92|93 => Pixel_t'(X"a",X"6",X"4"), 95 => Pixel_t'(X"a",X"a",X"b"), 43|91 => Pixel_t'(X"b",X"6",X"4"), 99 => Pixel_t'(X"d",X"d",X"f"), 96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    66 => (56 => Pixel_t'(X"4",X"3",X"2"), 26 => Pixel_t'(X"4",X"4",X"3"), 55|84 => Pixel_t'(X"5",X"3",X"2"), 57 => Pixel_t'(X"5",X"4",X"2"), 83 => Pixel_t'(X"5",X"4",X"3"), 58 => Pixel_t'(X"5",X"5",X"3"), 59|82 => Pixel_t'(X"5",X"6",X"4"), 85 => Pixel_t'(X"6",X"3",X"2"), 54 => Pixel_t'(X"6",X"4",X"2"), 94 => Pixel_t'(X"6",X"4",X"3"), 60|61 => Pixel_t'(X"6",X"7",X"4"), 81 => Pixel_t'(X"6",X"7",X"5"), 62|63|80 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24 => Pixel_t'(X"6",X"9",X"4"), 0|25|66|67|68|69|70|71|72|73|74|75|76|77 => Pixel_t'(X"6",X"9",X"5"), 53 => Pixel_t'(X"7",X"4",X"3"), 64|65|78|79 => Pixel_t'(X"7",X"9",X"5"), 27|52|86 => Pixel_t'(X"8",X"5",X"3"), 51|87 => Pixel_t'(X"9",X"6",X"4"), 30|44|91 => Pixel_t'(X"a",X"6",X"3"), 28|29|31|32|33|34|35|36|37|38|39|40|41|42|43|45|46|47|48|49|50|88|89|90|92|93 => Pixel_t'(X"a",X"6",X"4"), 95 => Pixel_t'(X"a",X"a",X"b"), 97|98|99 => Pixel_t'(X"d",X"d",X"f"), 96 => Pixel_t'(X"d",X"e",X"f")),
    67 => (63|80 => Pixel_t'(X"4",X"3",X"2"), 64|79 => Pixel_t'(X"4",X"4",X"2"), 26|61|62|81 => Pixel_t'(X"5",X"3",X"2"), 94 => Pixel_t'(X"5",X"4",X"4"), 65|66|78 => Pixel_t'(X"5",X"5",X"3"), 77 => Pixel_t'(X"5",X"5",X"4"), 67|68 => Pixel_t'(X"5",X"6",X"4"), 60 => Pixel_t'(X"6",X"4",X"3"), 76 => Pixel_t'(X"6",X"6",X"4"), 25|69|70|75 => Pixel_t'(X"6",X"7",X"4"), 71|72|73|74 => Pixel_t'(X"6",X"7",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 0|24 => Pixel_t'(X"6",X"9",X"5"), 59|82 => Pixel_t'(X"7",X"4",X"3"), 58 => Pixel_t'(X"8",X"4",X"3"), 83 => Pixel_t'(X"8",X"5",X"3"), 57 => Pixel_t'(X"9",X"5",X"3"), 33|56|84|93 => Pixel_t'(X"9",X"6",X"4"), 43|44|47|48|49|50|91 => Pixel_t'(X"a",X"6",X"3"), 27|28|29|30|31|32|34|35|36|37|38|39|40|41|42|45|46|51|52|53|54|55|85|86|87|88|89|90|92 => Pixel_t'(X"a",X"6",X"4"), 95 => Pixel_t'(X"d",X"c",X"d"), 97|98|99 => Pixel_t'(X"d",X"d",X"f"), 96 => Pixel_t'(X"d",X"e",X"f")),
    68 => (93 => Pixel_t'(X"5",X"3",X"3"), 25 => Pixel_t'(X"5",X"5",X"3"), 33|34|35|36|37 => Pixel_t'(X"6",X"2",X"2"), 32|38|70|71|72|74|75 => Pixel_t'(X"6",X"3",X"2"), 68|69|73 => Pixel_t'(X"6",X"4",X"2"), 76 => Pixel_t'(X"6",X"4",X"3"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 0|24 => Pixel_t'(X"6",X"9",X"5"), 39 => Pixel_t'(X"7",X"3",X"3"), 67 => Pixel_t'(X"7",X"4",X"2"), 66|77 => Pixel_t'(X"7",X"4",X"3"), 78 => Pixel_t'(X"8",X"4",X"3"), 40 => Pixel_t'(X"8",X"4",X"4"), 26|64|65|79 => Pixel_t'(X"8",X"5",X"3"), 63 => Pixel_t'(X"9",X"5",X"3"), 41 => Pixel_t'(X"9",X"5",X"4"), 80 => Pixel_t'(X"9",X"6",X"4"), 92 => Pixel_t'(X"9",X"6",X"5"), 94 => Pixel_t'(X"9",X"9",X"a"), 31 => Pixel_t'(X"a",X"5",X"3"), 50|51|52|53|54|56 => Pixel_t'(X"a",X"6",X"3"), 27|28|29|30|43|44|45|46|47|48|49|55|60|61|62|81|82|83|84|85|86|87|88|90|91 => Pixel_t'(X"a",X"6",X"4"), 42 => Pixel_t'(X"a",X"6",X"5"), 57 => Pixel_t'(X"b",X"6",X"3"), 58|59|89 => Pixel_t'(X"b",X"6",X"4"), 96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 95 => Pixel_t'(X"e",X"e",X"f")),
    69 => (92 => Pixel_t'(X"5",X"3",X"3"), 25 => Pixel_t'(X"5",X"4",X"3"), 41|42|43 => Pixel_t'(X"6",X"3",X"2"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23 => Pixel_t'(X"6",X"9",X"4"), 0|24 => Pixel_t'(X"6",X"9",X"5"), 40 => Pixel_t'(X"7",X"3",X"2"), 44 => Pixel_t'(X"7",X"4",X"3"), 39 => Pixel_t'(X"8",X"4",X"3"), 91 => Pixel_t'(X"8",X"5",X"4"), 38 => Pixel_t'(X"9",X"5",X"3"), 45 => Pixel_t'(X"9",X"5",X"4"), 26|33|35|36|37 => Pixel_t'(X"9",X"6",X"4"), 46 => Pixel_t'(X"9",X"6",X"5"), 93 => Pixel_t'(X"9",X"9",X"9"), 54|59|62|80|81 => Pixel_t'(X"a",X"6",X"3"), 27|28|29|30|31|32|34|48|49|50|51|52|53|55|56|57|58|60|61|63|64|65|66|68|69|70|71|72|73|74|75|76|78|82|83|84|85|86|87|89|90 => Pixel_t'(X"a",X"6",X"4"), 47 => Pixel_t'(X"a",X"6",X"5"), 79|88 => Pixel_t'(X"b",X"6",X"3"), 67|77 => Pixel_t'(X"b",X"6",X"4"), 95|96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 94 => Pixel_t'(X"e",X"e",X"f")),
    70 => (25 => Pixel_t'(X"5",X"4",X"2"), 91 => Pixel_t'(X"5",X"4",X"4"), 45|46|47 => Pixel_t'(X"6",X"3",X"2"), 90 => Pixel_t'(X"6",X"4",X"4"), 24 => Pixel_t'(X"6",X"8",X"5"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|23 => Pixel_t'(X"6",X"9",X"4"), 0|20|21|22 => Pixel_t'(X"6",X"9",X"5"), 44 => Pixel_t'(X"7",X"3",X"2"), 48 => Pixel_t'(X"7",X"3",X"3"), 43|49 => Pixel_t'(X"8",X"4",X"3"), 50 => Pixel_t'(X"9",X"5",X"4"), 42|51 => Pixel_t'(X"9",X"6",X"4"), 89 => Pixel_t'(X"9",X"6",X"5"), 32|78|79 => Pixel_t'(X"a",X"6",X"3"), 26|27|28|29|30|31|33|34|35|38|40|41|52|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|80|81|82|83|84|85|86|87 => Pixel_t'(X"a",X"6",X"4"), 53|88 => Pixel_t'(X"a",X"6",X"5"), 92 => Pixel_t'(X"a",X"a",X"b"), 36|37|39 => Pixel_t'(X"b",X"6",X"4"), 94|95|96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 93 => Pixel_t'(X"d",X"e",X"f")),
    71 => (89 => Pixel_t'(X"5",X"2",X"2"), 25 => Pixel_t'(X"5",X"4",X"2"), 90 => Pixel_t'(X"5",X"4",X"5"), 50|51 => Pixel_t'(X"6",X"2",X"2"), 52 => Pixel_t'(X"6",X"3",X"2"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|23 => Pixel_t'(X"6",X"9",X"4"), 0|20|21|22|24 => Pixel_t'(X"6",X"9",X"5"), 49|53 => Pixel_t'(X"7",X"3",X"2"), 54|87|88 => Pixel_t'(X"7",X"4",X"3"), 48 => Pixel_t'(X"8",X"4",X"3"), 55|86 => Pixel_t'(X"8",X"5",X"4"), 47|56|85 => Pixel_t'(X"9",X"5",X"4"), 57|84 => Pixel_t'(X"9",X"6",X"4"), 58 => Pixel_t'(X"9",X"6",X"5"), 29 => Pixel_t'(X"a",X"6",X"3"), 26|27|28|30|31|32|33|34|35|36|38|39|40|41|42|43|44|45|46|60|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|83 => Pixel_t'(X"a",X"6",X"4"), 59 => Pixel_t'(X"a",X"6",X"5"), 37 => Pixel_t'(X"b",X"6",X"4"), 91 => Pixel_t'(X"c",X"c",X"d"), 95 => Pixel_t'(X"d",X"d",X"e"), 94|96|97|98|99 => Pixel_t'(X"d",X"d",X"f"), 93 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    72 => (25 => Pixel_t'(X"5",X"5",X"3"), 57|84 => Pixel_t'(X"6",X"2",X"2"), 56|58|59|82|83|85 => Pixel_t'(X"6",X"3",X"2"), 1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|22|23 => Pixel_t'(X"6",X"9",X"4"), 0|20|21|24 => Pixel_t'(X"6",X"9",X"5"), 55|86 => Pixel_t'(X"7",X"3",X"2"), 60|81 => Pixel_t'(X"7",X"3",X"3"), 54 => Pixel_t'(X"7",X"4",X"2"), 61|62|63|78|79|80|87|89 => Pixel_t'(X"7",X"4",X"3"), 26 => Pixel_t'(X"7",X"5",X"3"), 90 => Pixel_t'(X"7",X"6",X"6"), 64|77 => Pixel_t'(X"8",X"4",X"3"), 53|65|66|76|88 => Pixel_t'(X"8",X"5",X"3"), 67|68|69|70|71|72|73|74|75 => Pixel_t'(X"8",X"5",X"4"), 52 => Pixel_t'(X"9",X"5",X"3"), 42|43|44 => Pixel_t'(X"a",X"6",X"3"), 28|29|30|31|32|33|34|35|36|37|38|39|40|41|45|46|47|48|49|50|51 => Pixel_t'(X"a",X"6",X"4"), 27 => Pixel_t'(X"a",X"6",X"5"), 92|93|94|95|96|97|99 => Pixel_t'(X"d",X"d",X"f"), 98 => Pixel_t'(X"d",X"e",X"f"), 91 => Pixel_t'(X"e",X"e",X"f")),
    73 => (26 => Pixel_t'(X"4",X"4",X"2"), 67|68|69|70|71|72|73|74 => Pixel_t'(X"6",X"3",X"2"), 90 => Pixel_t'(X"6",X"4",X"3"), 21 => Pixel_t'(X"6",X"8",X"4"), 25 => Pixel_t'(X"6",X"8",X"5"), 1|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|23|24 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|20|22 => Pixel_t'(X"6",X"9",X"5"), 65|66|75|76 => Pixel_t'(X"7",X"3",X"2"), 64|77|78 => Pixel_t'(X"7",X"4",X"2"), 27 => Pixel_t'(X"7",X"5",X"4"), 63 => Pixel_t'(X"8",X"4",X"2"), 61|62|79|80 => Pixel_t'(X"8",X"4",X"3"), 59|60|81 => Pixel_t'(X"9",X"5",X"3"), 58|82|83 => Pixel_t'(X"9",X"5",X"4"), 29|30 => Pixel_t'(X"9",X"6",X"4"), 28 => Pixel_t'(X"9",X"6",X"5"), 44 => Pixel_t'(X"a",X"6",X"3"), 31|37|38|39|40|41|42|43|47|48|49|50|51|52|53|54|55|56|57|84|85|86|87|88|89 => Pixel_t'(X"a",X"6",X"4"), 32|33|34|35|36 => Pixel_t'(X"a",X"6",X"5"), 45 => Pixel_t'(X"b",X"6",X"3"), 46 => Pixel_t'(X"b",X"6",X"4"), 91 => Pixel_t'(X"c",X"c",X"d"), 94|95|96|99 => Pixel_t'(X"d",X"d",X"f"), 92|93|97|98 => Pixel_t'(X"d",X"e",X"f")),
    74 => (28 => Pixel_t'(X"3",X"3",X"2"), 27 => Pixel_t'(X"3",X"4",X"2"), 21 => Pixel_t'(X"3",X"6",X"2"), 32|33|34|35|36 => Pixel_t'(X"4",X"3",X"2"), 29|30|31|37 => Pixel_t'(X"4",X"4",X"2"), 38 => Pixel_t'(X"5",X"4",X"3"), 90 => Pixel_t'(X"6",X"4",X"3"), 39 => Pixel_t'(X"6",X"5",X"3"), 22|26 => Pixel_t'(X"6",X"8",X"5"), 1|8|9|10|11|12|13|14|15|16|17|18|19|23|24 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|7|20|25 => Pixel_t'(X"6",X"9",X"5"), 40 => Pixel_t'(X"7",X"5",X"4"), 41|42 => Pixel_t'(X"9",X"6",X"4"), 47|48|49|85|86|87 => Pixel_t'(X"a",X"6",X"3"), 43|44|45|46|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|74|75|76|77|78|79|80|81|82|83|84|88|89 => Pixel_t'(X"a",X"6",X"4"), 91 => Pixel_t'(X"a",X"a",X"b"), 73 => Pixel_t'(X"b",X"6",X"4"), 93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    75 => (41|42 => Pixel_t'(X"4",X"4",X"2"), 40 => Pixel_t'(X"4",X"5",X"2"), 21|39 => Pixel_t'(X"4",X"6",X"3"), 22 => Pixel_t'(X"4",X"7",X"4"), 43 => Pixel_t'(X"5",X"4",X"2"), 90 => Pixel_t'(X"5",X"4",X"4"), 38 => Pixel_t'(X"5",X"6",X"4"), 37 => Pixel_t'(X"5",X"7",X"4"), 28|33|34|35|36 => Pixel_t'(X"5",X"8",X"4"), 44 => Pixel_t'(X"6",X"4",X"3"), 29|30|31|32 => Pixel_t'(X"6",X"8",X"4"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|24|25 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|20|23|26|27 => Pixel_t'(X"6",X"9",X"5"), 45 => Pixel_t'(X"8",X"5",X"4"), 46 => Pixel_t'(X"9",X"6",X"4"), 59|60|83|87 => Pixel_t'(X"a",X"6",X"3"), 48|49|50|51|52|54|55|56|57|58|61|62|63|64|65|66|67|68|69|70|71|72|73|74|75|76|77|78|79|80|81|82|84|85|86|88 => Pixel_t'(X"a",X"6",X"4"), 47|89 => Pixel_t'(X"a",X"6",X"5"), 53 => Pixel_t'(X"b",X"6",X"4"), 91 => Pixel_t'(X"c",X"c",X"d"), 93|99 => Pixel_t'(X"d",X"d",X"f"), 94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 92 => Pixel_t'(X"e",X"e",X"f")),
    76 => (22 => Pixel_t'(X"3",X"5",X"2"), 45|46 => Pixel_t'(X"4",X"4",X"2"), 44 => Pixel_t'(X"4",X"6",X"3"), 47 => Pixel_t'(X"5",X"4",X"2"), 43 => Pixel_t'(X"5",X"7",X"4"), 48 => Pixel_t'(X"6",X"4",X"3"), 90 => Pixel_t'(X"6",X"6",X"6"), 21|23|42 => Pixel_t'(X"6",X"8",X"5"), 1|7|8|9|10|11|12|13|14|15|16|17|18|19|25|26|27|28|29 => Pixel_t'(X"6",X"9",X"4"), 0|2|3|4|5|6|20|24|30|31|32|33|34|35|36|37|38|39|40|41 => Pixel_t'(X"6",X"9",X"5"), 89 => Pixel_t'(X"7",X"4",X"4"), 49 => Pixel_t'(X"7",X"5",X"4"), 50 => Pixel_t'(X"8",X"6",X"5"), 59|60|61|63|71|86|87 => Pixel_t'(X"a",X"6",X"3"), 53|54|55|56|57|58|62|64|65|66|67|68|69|70|72|73|74|75|76|77|78|79|80|81|82|83|84|85|88 => Pixel_t'(X"a",X"6",X"4"), 51|52 => Pixel_t'(X"a",X"6",X"5"), 92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 91|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    77 => (50 => Pixel_t'(X"3",X"4",X"2"), 51 => Pixel_t'(X"4",X"4",X"2"), 89 => Pixel_t'(X"4",X"4",X"4"), 49 => Pixel_t'(X"4",X"5",X"2"), 22|23|48 => Pixel_t'(X"4",X"6",X"3"), 52 => Pixel_t'(X"5",X"4",X"3"), 47 => Pixel_t'(X"5",X"7",X"4"), 53 => Pixel_t'(X"6",X"4",X"3"), 0 => Pixel_t'(X"6",X"8",X"4"), 46 => Pixel_t'(X"6",X"8",X"5"), 5|6|7|8|9|10|11|12|13|14|15|16|17|20|27|28|29|30|31|32|33|34|35|36|37|42|43|44 => Pixel_t'(X"6",X"9",X"4"), 1|2|3|4|18|19|21|24|25|26|38|39|40|41|45 => Pixel_t'(X"6",X"9",X"5"), 88 => Pixel_t'(X"7",X"4",X"4"), 54 => Pixel_t'(X"7",X"5",X"4"), 55 => Pixel_t'(X"8",X"5",X"4"), 57 => Pixel_t'(X"9",X"6",X"4"), 56 => Pixel_t'(X"9",X"6",X"5"), 74|75|76|77|78|79|82 => Pixel_t'(X"a",X"6",X"3"), 58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73|80|81|84|85|86|87 => Pixel_t'(X"a",X"6",X"4"), 83 => Pixel_t'(X"b",X"6",X"4"), 90 => Pixel_t'(X"c",X"c",X"d"), 92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 91|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    78 => (55|56 => Pixel_t'(X"3",X"4",X"2"), 23 => Pixel_t'(X"3",X"5",X"2"), 24 => Pixel_t'(X"3",X"6",X"3"), 57|58 => Pixel_t'(X"4",X"4",X"2"), 54 => Pixel_t'(X"4",X"5",X"3"), 0 => Pixel_t'(X"4",X"5",X"4"), 53 => Pixel_t'(X"4",X"6",X"3"), 59|60|87 => Pixel_t'(X"5",X"4",X"3"), 88 => Pixel_t'(X"5",X"5",X"5"), 52 => Pixel_t'(X"5",X"7",X"4"), 51 => Pixel_t'(X"5",X"8",X"4"), 61 => Pixel_t'(X"6",X"4",X"3"), 62 => Pixel_t'(X"6",X"5",X"3"), 1|25 => Pixel_t'(X"6",X"8",X"5"), 5|6|7|8|9|10|11|12|13|14|15|16|17|21|28|30|31|32|33|34|35|36|37|41|42|43|44|45|46|47 => Pixel_t'(X"6",X"9",X"4"), 2|3|4|18|19|20|22|27|29|38|39|40|48|49|50 => Pixel_t'(X"6",X"9",X"5"), 63 => Pixel_t'(X"7",X"5",X"3"), 64 => Pixel_t'(X"7",X"5",X"4"), 26 => Pixel_t'(X"7",X"9",X"5"), 65|66|86 => Pixel_t'(X"8",X"5",X"4"), 67 => Pixel_t'(X"8",X"6",X"4"), 69|70|85 => Pixel_t'(X"9",X"6",X"4"), 68 => Pixel_t'(X"9",X"6",X"5"), 73|74|75|76|77|78|79|80|81|82|83 => Pixel_t'(X"a",X"6",X"4"), 71|72|84 => Pixel_t'(X"a",X"6",X"5"), 89 => Pixel_t'(X"b",X"b",X"c"), 91|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 90 => Pixel_t'(X"e",X"e",X"f")),
    79 => (66|67|68|69|70|71 => Pixel_t'(X"3",X"4",X"2"), 25|65 => Pixel_t'(X"3",X"5",X"2"), 72|73|74|75 => Pixel_t'(X"4",X"4",X"2"), 64 => Pixel_t'(X"4",X"5",X"2"), 63 => Pixel_t'(X"4",X"5",X"3"), 24|26|62 => Pixel_t'(X"4",X"6",X"3"), 1 => Pixel_t'(X"4",X"6",X"4"), 83 => Pixel_t'(X"5",X"3",X"3"), 76|77 => Pixel_t'(X"5",X"4",X"2"), 78|79|80|82 => Pixel_t'(X"5",X"4",X"3"), 84|85 => Pixel_t'(X"5",X"4",X"4"), 61 => Pixel_t'(X"5",X"6",X"3"), 60 => Pixel_t'(X"5",X"7",X"3"), 27|59 => Pixel_t'(X"5",X"7",X"4"), 58 => Pixel_t'(X"5",X"8",X"4"), 81 => Pixel_t'(X"6",X"4",X"3"), 86 => Pixel_t'(X"6",X"5",X"6"), 57 => Pixel_t'(X"6",X"8",X"4"), 28 => Pixel_t'(X"6",X"8",X"5"), 3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|20|21|22|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52 => Pixel_t'(X"6",X"9",X"4"), 2|18|19|23|29|53|54|55|56 => Pixel_t'(X"6",X"9",X"5"), 0 => Pixel_t'(X"9",X"9",X"9"), 87 => Pixel_t'(X"9",X"9",X"a"), 88 => Pixel_t'(X"d",X"d",X"e"), 90|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 91 => Pixel_t'(X"e",X"d",X"f"), 89 => Pixel_t'(X"e",X"e",X"f")),
    80 => (81 => Pixel_t'(X"2",X"2",X"2"), 27 => Pixel_t'(X"3",X"6",X"2"), 26|28 => Pixel_t'(X"4",X"7",X"3"), 80 => Pixel_t'(X"5",X"6",X"4"), 2|74|75|76|77|78|79 => Pixel_t'(X"5",X"7",X"4"), 72|73 => Pixel_t'(X"5",X"8",X"4"), 82 => Pixel_t'(X"6",X"6",X"7"), 1 => Pixel_t'(X"6",X"7",X"6"), 70|71 => Pixel_t'(X"6",X"8",X"4"), 25|69 => Pixel_t'(X"6",X"8",X"5"), 4|5|6|7|8|9|10|11|12|13|14|15|19|20|21|22|23|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|55|56|57|58|59|60 => Pixel_t'(X"6",X"9",X"4"), 3|16|17|18|24|29|30|54|61|62|63|64|65|66|67|68 => Pixel_t'(X"6",X"9",X"5"), 83 => Pixel_t'(X"b",X"a",X"c"), 84 => Pixel_t'(X"b",X"b",X"d"), 85 => Pixel_t'(X"d",X"c",X"e"), 0 => Pixel_t'(X"d",X"d",X"e"), 88|89|90|91|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 86|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 87 => Pixel_t'(X"e",X"e",X"f")),
    81 => (2 => Pixel_t'(X"2",X"3",X"2"), 80 => Pixel_t'(X"4",X"5",X"4"), 3 => Pixel_t'(X"5",X"7",X"4"), 6|7|8|9|10|11|12|19|20|21|22|23|24|25|28|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|54|55|56|59|60|61|64|65|66|67|68|69|70|71|72|74|75 => Pixel_t'(X"6",X"9",X"4"), 4|5|13|14|15|16|17|18|26|27|29|53|57|58|62|63|73|76|77 => Pixel_t'(X"6",X"9",X"5"), 81 => Pixel_t'(X"7",X"7",X"8"), 78|79 => Pixel_t'(X"7",X"9",X"5"), 1 => Pixel_t'(X"8",X"8",X"8"), 85|87|88|89|90|91|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 82|86|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 0|83|84 => Pixel_t'(X"e",X"e",X"f")),
    82 => (1 => Pixel_t'(X"2",X"3",X"6"), 4 => Pixel_t'(X"3",X"5",X"2"), 79 => Pixel_t'(X"4",X"5",X"3"), 3 => Pixel_t'(X"4",X"6",X"3"), 0 => Pixel_t'(X"5",X"5",X"a"), 2 => Pixel_t'(X"5",X"6",X"5"), 5 => Pixel_t'(X"5",X"7",X"4"), 78 => Pixel_t'(X"6",X"8",X"5"), 8|9|10|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|59|64|65|66|67|68|69|70|71|72|76 => Pixel_t'(X"6",X"9",X"4"), 6|7|11|12|13|14|15|16|17|18|56|57|58|60|61|62|63|73|74|75 => Pixel_t'(X"6",X"9",X"5"), 80 => Pixel_t'(X"7",X"8",X"8"), 77 => Pixel_t'(X"7",X"9",X"5"), 81|83|84|85|88|89|90|91|92|93|94|99 => Pixel_t'(X"d",X"d",X"f"), 86 => Pixel_t'(X"d",X"e",X"e"), 82|87|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    83 => (1 => Pixel_t'(X"1",X"3",X"b"), 2 => Pixel_t'(X"2",X"3",X"7"), 0 => Pixel_t'(X"2",X"3",X"d"), 78 => Pixel_t'(X"3",X"4",X"3"), 5 => Pixel_t'(X"3",X"5",X"2"), 6 => Pixel_t'(X"3",X"5",X"3"), 7 => Pixel_t'(X"5",X"8",X"4"), 4|77 => Pixel_t'(X"6",X"7",X"5"), 3 => Pixel_t'(X"6",X"7",X"6"), 10|11|12|13|14|15|16|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|62|63|64|65|69|70|71|72|73|74|75 => Pixel_t'(X"6",X"9",X"4"), 8|9|17|18|57|58|59|60|61|66|67|68 => Pixel_t'(X"6",X"9",X"5"), 76 => Pixel_t'(X"7",X"9",X"5"), 79 => Pixel_t'(X"8",X"9",X"9"), 81|82|83|84|90|91|92|93|99 => Pixel_t'(X"d",X"d",X"f"), 85|86|87|88|89|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 80 => Pixel_t'(X"e",X"e",X"f")),
    84 => (3 => Pixel_t'(X"1",X"3",X"7"), 2 => Pixel_t'(X"2",X"4",X"c"), 0|1 => Pixel_t'(X"2",X"4",X"f"), 7 => Pixel_t'(X"3",X"5",X"2"), 8 => Pixel_t'(X"3",X"6",X"3"), 77 => Pixel_t'(X"4",X"4",X"4"), 76 => Pixel_t'(X"4",X"5",X"4"), 4 => Pixel_t'(X"4",X"6",X"6"), 6|9 => Pixel_t'(X"5",X"7",X"4"), 13|14|15|16|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|44|45|46|47|48|49|50|51|52|53|54|55|61|62|63|64|69|70|71|72|73 => Pixel_t'(X"6",X"9",X"4"), 10|12|17|18|41|42|43|56|57|58|59|60|65|66|67|68 => Pixel_t'(X"6",X"9",X"5"), 75 => Pixel_t'(X"7",X"8",X"5"), 5 => Pixel_t'(X"7",X"8",X"6"), 11|74 => Pixel_t'(X"7",X"9",X"5"), 78 => Pixel_t'(X"a",X"b",X"b"), 80|81|82|83|84|90|91|92|93|99 => Pixel_t'(X"d",X"d",X"f"), 85|86|87|88|89|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 79 => Pixel_t'(X"e",X"e",X"f")),
    85 => (4 => Pixel_t'(X"1",X"3",X"9"), 3 => Pixel_t'(X"2",X"4",X"d"), 0|1|2 => Pixel_t'(X"2",X"4",X"f"), 75 => Pixel_t'(X"3",X"4",X"3"), 5 => Pixel_t'(X"3",X"4",X"6"), 9|10 => Pixel_t'(X"3",X"5",X"2"), 8|11 => Pixel_t'(X"5",X"7",X"4"), 74 => Pixel_t'(X"5",X"7",X"5"), 76 => Pixel_t'(X"6",X"7",X"7"), 12 => Pixel_t'(X"6",X"8",X"5"), 6 => Pixel_t'(X"6",X"8",X"6"), 16|17|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|44|45|46|47|48|49|50|51|52|53|54|55|62|63|64|69|70 => Pixel_t'(X"6",X"9",X"4"), 13|14|15|18|41|42|43|56|57|58|59|60|61|65|66|67|68|71|72 => Pixel_t'(X"6",X"9",X"5"), 7 => Pixel_t'(X"7",X"8",X"5"), 73 => Pixel_t'(X"7",X"9",X"5"), 77 => Pixel_t'(X"c",X"c",X"e"), 79|80|81|82|83|84|90|91|92|99 => Pixel_t'(X"d",X"d",X"f"), 85|86|87|88|89|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 78 => Pixel_t'(X"e",X"e",X"f")),
    86 => (6 => Pixel_t'(X"1",X"3",X"7"), 5 => Pixel_t'(X"1",X"3",X"c"), 4 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3 => Pixel_t'(X"2",X"4",X"f"), 12 => Pixel_t'(X"2",X"5",X"2"), 13 => Pixel_t'(X"3",X"6",X"3"), 73 => Pixel_t'(X"4",X"5",X"3"), 11 => Pixel_t'(X"4",X"6",X"3"), 7 => Pixel_t'(X"4",X"6",X"6"), 74 => Pixel_t'(X"5",X"5",X"5"), 10|14 => Pixel_t'(X"5",X"7",X"4"), 72 => Pixel_t'(X"6",X"7",X"5"), 15 => Pixel_t'(X"6",X"8",X"5"), 8 => Pixel_t'(X"6",X"8",X"6"), 20|21|22|23|24|25|28|29|30|31|32|33|34|35|36|37|38|39|40|41|44|45|46|47|48|49|50|51|52|53|54|55|62|63|67|68|69 => Pixel_t'(X"6",X"9",X"4"), 16|17|18|19|26|27|42|43|56|57|58|59|60|61|64|65|66|70 => Pixel_t'(X"6",X"9",X"5"), 9|71 => Pixel_t'(X"7",X"9",X"5"), 75 => Pixel_t'(X"a",X"a",X"b"), 78|79|80|81|82|83|84|99 => Pixel_t'(X"d",X"d",X"f"), 76|77|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")),
    87 => (7 => Pixel_t'(X"1",X"3",X"a"), 8 => Pixel_t'(X"2",X"3",X"6"), 6 => Pixel_t'(X"2",X"4",X"d"), 0|1|2|3|4|5 => Pixel_t'(X"2",X"4",X"f"), 71 => Pixel_t'(X"3",X"4",X"3"), 15 => Pixel_t'(X"3",X"5",X"2"), 16 => Pixel_t'(X"3",X"5",X"3"), 14 => Pixel_t'(X"3",X"6",X"2"), 17 => Pixel_t'(X"4",X"7",X"4"), 72 => Pixel_t'(X"5",X"5",X"5"), 13 => Pixel_t'(X"5",X"7",X"3"), 70 => Pixel_t'(X"5",X"7",X"5"), 9 => Pixel_t'(X"5",X"7",X"6"), 18 => Pixel_t'(X"5",X"8",X"4"), 12|19 => Pixel_t'(X"6",X"8",X"5"), 25|26|27|28|29|31|32|33|34|35|36|37|38|39|40|46|47|48|49|50|51|52|53|54|55|62|63|64|65 => Pixel_t'(X"6",X"9",X"4"), 20|21|22|23|24|30|41|42|43|44|45|56|57|58|59|60|61|66|67 => Pixel_t'(X"6",X"9",X"5"), 10 => Pixel_t'(X"6",X"9",X"6"), 11|68|69 => Pixel_t'(X"7",X"9",X"5"), 73 => Pixel_t'(X"a",X"a",X"a"), 74 => Pixel_t'(X"d",X"d",X"e"), 76|77|78|79|80|81|82|83|99 => Pixel_t'(X"d",X"d",X"f"), 84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 75 => Pixel_t'(X"e",X"e",X"f")),
    88 => (9 => Pixel_t'(X"1",X"3",X"9"), 8 => Pixel_t'(X"1",X"3",X"d"), 10 => Pixel_t'(X"2",X"4",X"6"), 0|1|2|3|4|5|6|7 => Pixel_t'(X"2",X"4",X"f"), 69 => Pixel_t'(X"3",X"4",X"3"), 18|19|20 => Pixel_t'(X"3",X"5",X"2"), 17 => Pixel_t'(X"3",X"6",X"3"), 21 => Pixel_t'(X"4",X"6",X"3"), 68 => Pixel_t'(X"4",X"6",X"4"), 70 => Pixel_t'(X"5",X"6",X"5"), 16 => Pixel_t'(X"5",X"7",X"3"), 22 => Pixel_t'(X"5",X"7",X"4"), 11 => Pixel_t'(X"5",X"7",X"6"), 23 => Pixel_t'(X"5",X"8",X"5"), 67 => Pixel_t'(X"6",X"7",X"5"), 15 => Pixel_t'(X"6",X"8",X"4"), 24 => Pixel_t'(X"6",X"8",X"5"), 29|33|34|35|36|37|38|39|46|47|48|49|50|51|52|53|54|55|59|60|61|62|63|64|65 => Pixel_t'(X"6",X"9",X"4"), 14|25|26|28|30|31|32|40|41|42|43|44|45|56|57|58 => Pixel_t'(X"6",X"9",X"5"), 13|27|66 => Pixel_t'(X"7",X"9",X"5"), 12 => Pixel_t'(X"7",X"9",X"6"), 71 => Pixel_t'(X"9",X"9",X"a"), 72 => Pixel_t'(X"d",X"d",X"e"), 74|75|76|77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 73 => Pixel_t'(X"e",X"e",X"f")),
    89 => (11 => Pixel_t'(X"1",X"2",X"9"), 10 => Pixel_t'(X"2",X"3",X"c"), 0|1|2|3|4|5|6|7|8|9 => Pixel_t'(X"2",X"4",X"f"), 12 => Pixel_t'(X"3",X"4",X"7"), 23|24|25 => Pixel_t'(X"3",X"5",X"2"), 26 => Pixel_t'(X"3",X"5",X"3"), 22 => Pixel_t'(X"3",X"6",X"2"), 66 => Pixel_t'(X"4",X"5",X"4"), 27 => Pixel_t'(X"4",X"6",X"3"), 21 => Pixel_t'(X"4",X"7",X"3"), 67 => Pixel_t'(X"5",X"5",X"5"), 28 => Pixel_t'(X"5",X"6",X"4"), 29 => Pixel_t'(X"5",X"7",X"4"), 13 => Pixel_t'(X"5",X"7",X"6"), 20 => Pixel_t'(X"5",X"8",X"4"), 19|30|31 => Pixel_t'(X"6",X"8",X"5"), 46|47|48|49|50|51|52|53|54|55 => Pixel_t'(X"6",X"9",X"4"), 14|17|18|32|33|34|35|36|37|38|39|40|41|42|43|44|45|56|57|58|59|60|61|62|63 => Pixel_t'(X"6",X"9",X"5"), 15|16|64 => Pixel_t'(X"7",X"9",X"5"), 65 => Pixel_t'(X"7",X"9",X"6"), 68 => Pixel_t'(X"8",X"8",X"9"), 69 => Pixel_t'(X"a",X"a",X"b"), 70 => Pixel_t'(X"d",X"d",X"e"), 73|74|76|77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 75|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 72 => Pixel_t'(X"e",X"d",X"f"), 71 => Pixel_t'(X"e",X"e",X"f")),
    90 => (13 => Pixel_t'(X"1",X"2",X"9"), 64 => Pixel_t'(X"2",X"3",X"4"), 65 => Pixel_t'(X"2",X"3",X"5"), 14 => Pixel_t'(X"2",X"3",X"7"), 12 => Pixel_t'(X"2",X"3",X"c"), 11 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10 => Pixel_t'(X"2",X"4",X"f"), 31 => Pixel_t'(X"2",X"5",X"2"), 29|30 => Pixel_t'(X"3",X"5",X"2"), 32|63 => Pixel_t'(X"3",X"5",X"3"), 33 => Pixel_t'(X"3",X"6",X"3"), 28|34|35|61|62 => Pixel_t'(X"4",X"6",X"3"), 36 => Pixel_t'(X"4",X"6",X"4"), 15 => Pixel_t'(X"4",X"6",X"6"), 27 => Pixel_t'(X"4",X"7",X"3"), 66 => Pixel_t'(X"5",X"6",X"7"), 37|38|60 => Pixel_t'(X"5",X"7",X"4"), 26|59 => Pixel_t'(X"5",X"8",X"4"), 25 => Pixel_t'(X"6",X"8",X"4"), 39|40|41|42|57|58 => Pixel_t'(X"6",X"8",X"5"), 16 => Pixel_t'(X"6",X"8",X"6"), 19|21 => Pixel_t'(X"6",X"9",X"4"), 17|18|20|22|23|24|43|47|48|49|50|51|52|53|54|55|56 => Pixel_t'(X"6",X"9",X"5"), 44|45|46 => Pixel_t'(X"7",X"9",X"5"), 67 => Pixel_t'(X"d",X"d",X"e"), 71|72|73|74|99 => Pixel_t'(X"d",X"d",X"f"), 70 => Pixel_t'(X"d",X"e",X"e"), 75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 68|69 => Pixel_t'(X"e",X"e",X"f")),
    91 => (64 => Pixel_t'(X"1",X"2",X"8"), 65 => Pixel_t'(X"1",X"2",X"9"), 16 => Pixel_t'(X"1",X"3",X"8"), 15 => Pixel_t'(X"1",X"3",X"9"), 14 => Pixel_t'(X"2",X"4",X"d"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'(X"2",X"4",X"f"), 58 => Pixel_t'(X"3",X"4",X"2"), 37|38|39|40|41|42|43|44|45|53|54|55|56|57|59|60 => Pixel_t'(X"3",X"5",X"2"), 46|47|48|52 => Pixel_t'(X"3",X"5",X"3"), 17 => Pixel_t'(X"3",X"5",X"6"), 50|51 => Pixel_t'(X"3",X"6",X"3"), 63 => Pixel_t'(X"4",X"5",X"6"), 35|36|49|61 => Pixel_t'(X"4",X"6",X"3"), 34|62 => Pixel_t'(X"5",X"7",X"4"), 18 => Pixel_t'(X"5",X"7",X"6"), 33 => Pixel_t'(X"5",X"8",X"4"), 66 => Pixel_t'(X"6",X"7",X"a"), 32 => Pixel_t'(X"6",X"8",X"4"), 19 => Pixel_t'(X"6",X"8",X"5"), 22|24|25|26|27|31 => Pixel_t'(X"6",X"9",X"4"), 20|21|23|28|29|30 => Pixel_t'(X"6",X"9",X"5"), 70|71|72|99 => Pixel_t'(X"d",X"d",X"f"), 68|69|73|74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 67 => Pixel_t'(X"e",X"e",X"f")),
    92 => (66 => Pixel_t'(X"1",X"2",X"9"), 18 => Pixel_t'(X"1",X"3",X"9"), 17 => Pixel_t'(X"1",X"3",X"c"), 64 => Pixel_t'(X"1",X"4",X"d"), 19 => Pixel_t'(X"2",X"3",X"7"), 63 => Pixel_t'(X"2",X"3",X"8"), 16|65 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15 => Pixel_t'(X"2",X"4",X"f"), 20 => Pixel_t'(X"3",X"4",X"6"), 21 => Pixel_t'(X"5",X"6",X"6"), 47|48|49|50|51 => Pixel_t'(X"5",X"7",X"4"), 44|45|46|52|53|54|55 => Pixel_t'(X"5",X"8",X"4"), 67 => Pixel_t'(X"6",X"6",X"a"), 22 => Pixel_t'(X"6",X"7",X"6"), 62 => Pixel_t'(X"6",X"7",X"7"), 43|56|57 => Pixel_t'(X"6",X"8",X"4"), 42 => Pixel_t'(X"6",X"8",X"5"), 23 => Pixel_t'(X"6",X"8",X"6"), 29|30|31|32|33|34|35|40|41 => Pixel_t'(X"6",X"9",X"4"), 24|25|26|27|28|36|37|38|39|58|59 => Pixel_t'(X"6",X"9",X"5"), 60 => Pixel_t'(X"7",X"9",X"5"), 61 => Pixel_t'(X"7",X"9",X"6"), 68|70|71|72|73|99 => Pixel_t'(X"d",X"d",X"f"), 74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 69 => Pixel_t'(X"e",X"e",X"f")),
    93 => (67 => Pixel_t'(X"1",X"2",X"a"), 22 => Pixel_t'(X"1",X"3",X"8"), 62 => Pixel_t'(X"1",X"3",X"9"), 21 => Pixel_t'(X"1",X"3",X"a"), 20 => Pixel_t'(X"1",X"3",X"c"), 63 => Pixel_t'(X"1",X"3",X"d"), 23 => Pixel_t'(X"2",X"3",X"7"), 19|66 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|64|65 => Pixel_t'(X"2",X"4",X"f"), 24|61 => Pixel_t'(X"3",X"4",X"6"), 25 => Pixel_t'(X"3",X"5",X"6"), 68 => Pixel_t'(X"4",X"4",X"9"), 26 => Pixel_t'(X"4",X"6",X"6"), 27 => Pixel_t'(X"5",X"6",X"6"), 60 => Pixel_t'(X"5",X"7",X"6"), 28 => Pixel_t'(X"6",X"7",X"6"), 29|30|31|59 => Pixel_t'(X"6",X"8",X"6"), 38|39|40|41 => Pixel_t'(X"6",X"9",X"4"), 36|37|42|43|44|45|46|47|48|49|50|51|52|54|55|56|58 => Pixel_t'(X"6",X"9",X"5"), 32|33|34|35|53|57 => Pixel_t'(X"7",X"9",X"5"), 69 => Pixel_t'(X"b",X"b",X"d"), 72|73|99 => Pixel_t'(X"d",X"d",X"f"), 74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 71 => Pixel_t'(X"e",X"d",X"f"), 70 => Pixel_t'(X"e",X"e",X"f")),
    94 => (60 => Pixel_t'(X"1",X"2",X"a"), 29 => Pixel_t'(X"1",X"3",X"8"), 28 => Pixel_t'(X"1",X"3",X"9"), 26|27 => Pixel_t'(X"1",X"3",X"a"), 25 => Pixel_t'(X"1",X"3",X"b"), 24|61|68 => Pixel_t'(X"1",X"3",X"c"), 31 => Pixel_t'(X"2",X"3",X"7"), 30|59 => Pixel_t'(X"2",X"3",X"8"), 69 => Pixel_t'(X"2",X"3",X"9"), 22|23|62 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|63|64|65|66|67 => Pixel_t'(X"2",X"4",X"f"), 33 => Pixel_t'(X"3",X"4",X"6"), 32|58 => Pixel_t'(X"3",X"4",X"7"), 34|35|57 => Pixel_t'(X"4",X"5",X"6"), 36|56 => Pixel_t'(X"5",X"6",X"6"), 37|55 => Pixel_t'(X"5",X"7",X"6"), 38|39|54 => Pixel_t'(X"6",X"7",X"6"), 40|41|42|43|44|51|52|53 => Pixel_t'(X"6",X"8",X"6"), 45|46|47|48|49|50 => Pixel_t'(X"6",X"9",X"6"), 70 => Pixel_t'(X"8",X"8",X"b"), 71|73|99 => Pixel_t'(X"d",X"d",X"f"), 74|75|76|77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 72 => Pixel_t'(X"e",X"e",X"f")),
    95 => (38|55 => Pixel_t'(X"1",X"2",X"9"), 36|37|70 => Pixel_t'(X"1",X"2",X"a"), 39|54 => Pixel_t'(X"1",X"3",X"9"), 56 => Pixel_t'(X"1",X"3",X"a"), 34|35 => Pixel_t'(X"1",X"3",X"b"), 33|57 => Pixel_t'(X"1",X"3",X"c"), 32|58 => Pixel_t'(X"1",X"3",X"d"), 43|44|51 => Pixel_t'(X"2",X"3",X"7"), 40|41|42|52|53 => Pixel_t'(X"2",X"3",X"8"), 45|48|49|50 => Pixel_t'(X"2",X"4",X"7"), 46|47 => Pixel_t'(X"2",X"4",X"8"), 31|69 => Pixel_t'(X"2",X"4",X"d"), 29|30|59 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|60|61|62|63|64|65|66|67|68 => Pixel_t'(X"2",X"4",X"f"), 71 => Pixel_t'(X"5",X"5",X"9"), 72 => Pixel_t'(X"c",X"c",X"e"), 74|75|76|99 => Pixel_t'(X"d",X"d",X"f"), 77|78|79|80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 73 => Pixel_t'(X"e",X"e",X"f")),
    96 => (71 => Pixel_t'(X"1",X"3",X"b"), 46|47 => Pixel_t'(X"1",X"4",X"d"), 45 => Pixel_t'(X"1",X"4",X"e"), 72 => Pixel_t'(X"2",X"3",X"8"), 48|49 => Pixel_t'(X"2",X"4",X"d"), 39|40|41|42|43|44|50|51|52|53|54 => Pixel_t'(X"2",X"4",X"e"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70 => Pixel_t'(X"2",X"4",X"f"), 73 => Pixel_t'(X"a",X"a",X"d"), 75|76|77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 74 => Pixel_t'(X"e",X"e",X"f")),
    97 => (72 => Pixel_t'(X"1",X"3",X"c"), 73 => Pixel_t'(X"2",X"2",X"9"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71 => Pixel_t'(X"2",X"4",X"f"), 74 => Pixel_t'(X"a",X"a",X"c"), 76|77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 75 => Pixel_t'(X"e",X"e",X"f")),
    98 => (73 => Pixel_t'(X"1",X"3",X"d"), 74 => Pixel_t'(X"2",X"3",X"8"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72 => Pixel_t'(X"2",X"4",X"f"), 75 => Pixel_t'(X"b",X"a",X"d"), 77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f"), 76 => Pixel_t'(X"e",X"e",X"f")),
    99 => (74 => Pixel_t'(X"2",X"3",X"c"), 0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'(X"2",X"4",X"f"), 75 => Pixel_t'(X"3",X"3",X"8"), 76 => Pixel_t'(X"c",X"d",X"e"), 77|78|79|99 => Pixel_t'(X"d",X"d",X"f"), 80|81|82|83|84|85|86|87|88|89|90|91|92|93|94|95|96|97|98 => Pixel_t'(X"d",X"e",X"f")));


end package;