(0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
2 => (0|1|2|3|4|5|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 6|36|55|56 => Pixel_t'("01","01","01"), 11|12|13|14|15|31|32|33|34 => Pixel_t'("01","10","10"), 7|8|9|10|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|35 => Pixel_t'("10","10","10")),
3 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 53 => Pixel_t'("00","01","01"), 21|22|29 => Pixel_t'("01","01","01"), 19|20|23|24|25|26|28 => Pixel_t'("01","01","10"), 17|18|27 => Pixel_t'("01","10","10"), 1|2|3|4|5|12|13|14|15|16|30|31|32|33|34|35|36|54|55|57 => Pixel_t'("10","10","10"), 6 => Pixel_t'("10","10","11"), 56 => Pixel_t'("10","11","10"), 7|8 => Pixel_t'("10","11","11"), 9|10|11 => Pixel_t'("11","11","11")),
4 => (0|1|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|32|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","00","01"), 11|31|33|36|52 => Pixel_t'("01","01","01"), 5 => Pixel_t'("01","01","10"), 2|30 => Pixel_t'("01","10","10"), 3|4|6|7|34|35|53|54|55|56|57|58 => Pixel_t'("10","10","10"), 8 => Pixel_t'("10","10","11"), 9|10 => Pixel_t'("11","11","11")),
5 => (0|1|18|19|20|21|22|23|24|25|26|27|36|37|38|39|40|41|42|43|44|45|46|47|48|49|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 17 => Pixel_t'("00","00","01"), 16|28 => Pixel_t'("00","01","01"), 2|3|11|12|13|14|15|29|30|31|32|50|61 => Pixel_t'("01","01","01"), 51|60 => Pixel_t'("01","10","10"), 4|5|6|7|8|9|10|33|34|35|52|53|54|55|56|57|58|59 => Pixel_t'("10","10","10")),
6 => (0|1|2|5|6|7|8|9|10|36|37|44|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 3|4|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|39|40|41|43|45|46|47|65|66|67 => Pixel_t'("01","01","01"), 38|42|48|51|52|53|54|55|56|57|58|64 => Pixel_t'("01","10","10"), 49|50|59|60|61|62|63 => Pixel_t'("10","10","10")),
7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|19|28|29|30|31|32|33|34|35|36|37|73 => Pixel_t'("00","00","00"), 26|43|44 => Pixel_t'("00","01","01"), 18|20|21|22|23|24|25|27|38|41|42|45|46|47|48|49|50|51|52|53|54|55|56|57 => Pixel_t'("01","01","01"), 58|72 => Pixel_t'("01","01","10"), 39|40|59|60|61|62|63|64|65|66|67|68|69|70|71 => Pixel_t'("10","10","10")),
8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|26|27|28|29|30|31|32|33|34|35|36|37|38|49|50|51|52|64|67|68|73 => Pixel_t'("00","00","00"), 21|65|70 => Pixel_t'("00","00","01"), 53|66|69 => Pixel_t'("00","01","01"), 22|23|24|25|42|43|44|45|46|47|48|54|55|56|57|58|59|60|61|62|63|71|72 => Pixel_t'("01","01","01"), 39 => Pixel_t'("01","10","01"), 40|41 => Pixel_t'("10","10","10")),
9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|27|28|29|30|31|32|33|34|35|36|37|48|49|50|51|52|53|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 58 => Pixel_t'("00","01","01"), 24|25|26|47|54|57 => Pixel_t'("01","01","01"), 38|39|42|44|45|46|55|56 => Pixel_t'("10","10","10"), 43 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|28|29|30|31|32|33|34|35|36|47|48|49|50|51|52|53|54|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 25|26|27|46|57|58 => Pixel_t'("01","01","01"), 37|42|45|55|56 => Pixel_t'("10","10","10"), 38|44 => Pixel_t'("10","10","11"), 39|43 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|29|30|31|32|33|34|35|45|46|47|48|49|50|51|52|53|54|55|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 26 => Pixel_t'("00","01","01"), 27|28|56 => Pixel_t'("01","01","01"), 36|38|39|42|43|44 => Pixel_t'("10","10","10"), 37 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|31|32|33|34|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 30|35 => Pixel_t'("00","01","01"), 28|29 => Pixel_t'("01","01","01"), 36|37|38|39|40|42|43 => Pixel_t'("10","10","10"), 41 => Pixel_t'("10","11","11")),
13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|32|33|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29|30|31|34 => Pixel_t'("01","01","01"), 35|36 => Pixel_t'("01","10","10"), 37|38|39|40|41|42|43 => Pixel_t'("10","10","10")),
14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 30|31|32|33|34|35|36|37|38|39|40 => Pixel_t'("01","01","01"), 41|42 => Pixel_t'("01","10","10"), 43 => Pixel_t'("10","10","10")),
15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|30|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","01","01"), 21|22|23|24|31|32|44 => Pixel_t'("01","01","01"), 25|28|43 => Pixel_t'("01","10","10"), 26|27|33|34|35|36|37|38|39|40|41|42 => Pixel_t'("10","10","10")),
16 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 20|45 => Pixel_t'("01","01","01"), 43|44 => Pixel_t'("01","10","10"), 29|42 => Pixel_t'("10","10","10"), 21 => Pixel_t'("10","11","10"), 22|23|24|25|26|27|28|30|31|35|36|41 => Pixel_t'("10","11","11"), 32|33|34|37|38|39|40 => Pixel_t'("11","11","11")),
17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 45 => Pixel_t'("01","10","10"), 20|34|35|44 => Pixel_t'("10","10","10"), 22|23|24|25|26|27|28|29|30|31|32|33|36|37|38|43 => Pixel_t'("10","11","11"), 21|39|40|41|42 => Pixel_t'("11","11","11")),
18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 45 => Pixel_t'("01","01","01"), 20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|44 => Pixel_t'("10","10","10"), 40 => Pixel_t'("11","10","10"), 41|42|43 => Pixel_t'("11","11","11")),
19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 23|24|44|45 => Pixel_t'("01","01","01"), 27 => Pixel_t'("01","10","01"), 25|26|28|29|30|31|43 => Pixel_t'("01","10","10"), 32|33|34|35|36|37|38|39|40|42 => Pixel_t'("10","10","10"), 41 => Pixel_t'("11","11","11")),
20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 44 => Pixel_t'("00","01","01"), 27|28|29|30|31|32|33|34|35|36|41|42|43 => Pixel_t'("01","01","01"), 38 => Pixel_t'("01","01","10"), 37|39 => Pixel_t'("01","10","10"), 40 => Pixel_t'("10","10","10")),
21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 34|35|36|37|38|40|41|42|43|44 => Pixel_t'("01","01","01"), 39 => Pixel_t'("01","01","10")),
22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 42 => Pixel_t'("00","00","01"), 41 => Pixel_t'("00","01","01"), 38|39|40|43 => Pixel_t'("01","01","01")),
23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")));