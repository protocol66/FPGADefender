library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.my_data_types.all;

package bitmaps is
    constant BACKGROUND : Pixel_t := BLACK;
    constant MAIN_CLK_FREQ : integer := 50000000;

    constant screen_HEIGHT : positive := 479;
    constant screen_WIDTH : positive := 639;

    constant pepe_sizeX : positive := 100;
    constant pepe_sizeY : positive := 100;

    constant line_sizeX : positive := screen_WIDTH;
    constant line_sizeY : positive := 2;

    constant ship_sizeX : positive := 74;
    constant ship_sizeY : positive := 25;
    
    constant laser_sizeX : positive := 20;
    constant laser_sizeY : positive := 1;

    constant score_sizeX : positive := 15;
    constant score_sizeY : positive := 25;
    constant score_space_size :positive := 5;
    constant score_board_sizeX : positive := (score_sizeX + score_space_size)*5 + score_sizeY;
    constant score_board_sizeY : positive := score_sizeY;

    constant alien1_sizeX : positive := 40;
    constant alien1_sizeY : positive := 30;

    constant alien2_sizeX : positive := 30;
    constant alien2_sizeY : positive := 20;

    constant alien3_sizeX : positive := 10;
    constant alien3_sizeY : positive := 10;

    constant asteroid_sizeX : positive := 40;
    constant asteroid_sizeY : positive := 40;

    constant H_LINE : bit_map_t (0 to line_sizeY-1, 0 to line_sizeX-1) := (others => (others => WHITE));
    -- constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) := (others => (others => TEAL));
    constant LASER : bit_map_t (0 to laser_sizeY-1, 0 to laser_sizeX-1) := (others => (others => GREEN));
    -- constant ALIEN_1 : bit_map_t (0 to alien1_sizeY-1, 0 to alien1_sizeX-1) := (others => (others => YELLOW));
    -- constant ALIEN_2 : bit_map_t (0 to alien2_sizeY-1, 0 to alien2_sizeX-1) := (others => (others => RED)); 
    -- constant ALIEN_3 : bit_map_t (0 to alien3_sizeY-1, 0 to alien3_sizeX-1) := (others => (others => BLUE));  
    -- constant ASTEROID : bit_map_t (0 to asteroid_sizeY-1, 0 to asteroid_sizeX-1) := (others => (others => PURPLE)); 
    constant SATELLITE : bit_map_t (0 to asteroid_sizeY-1, 0 to asteroid_sizeX-1) := (others => (others => GREEN)); 

    constant fx1 : Sound_FX_t := (18, (550, 404, 315, 494, 182, 260, 455, 387, 340, 550, 404, 315, 494, 182, 260, 455, 387, 340, others => 0));
    constant fx2 : Sound_FX_t := (10, (300, 350, 500, 700, 990, 970, 1050, 1010, 950, 800, 770, 640, 500, 350, 355, others => 0));
    constant fx3 : Sound_FX_t := (6,  (500, 790, 950, 1300, 1710, 1650, 1300, 800, 700, others=> 0));
    constant fx4 : Sound_FX_t := (60, (1300, 1650, 1660, 1510, 1309, 1158, 1007, 855, others=> 0));
    constant fx5 : Sound_FX_t := (25, (300, 210, 310, 170, 250, 210, 310, 120, 220, 170, 160, 90, 290, 230, 140, 320, 200, 100, 250, 290, others => 0));
    constant fx6 : Sound_FX_t := (15, (700, 702, 698, 701, 699, 700, 250, 251, 249, 252, 248, 130, 131, 129, 132, 128, 130, 130, others=>0));

    -- constant score_9 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    -- constant score_8 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    -- constant score_7 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    -- constant score_6 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    -- constant score_5 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => PURPLE));
    -- constant score_4 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => YELLOW));
    -- constant score_3 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => RED));
    -- constant score_2 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BLUE));
    -- constant score_1 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => GREEN));
    -- constant score_0 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => TEAL));
    constant score_blank : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := (others => (others => BACKGROUND));
    
    -- DONT USE THIS... adds 30+ min to compile time...
    constant SHIP : bit_map_t (0 to ship_sizeY-1, 0 to ship_sizeX-1) :=
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
        1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
        2 => (0|1|2|3|4|5|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 6|36|55|56 => Pixel_t'("01","01","01"), 11|12|13|14|15|31|32|33|34 => Pixel_t'("01","10","10"), 7|8|9|10|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|35 => Pixel_t'("10","10","10")),
        3 => (0|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 53 => Pixel_t'("00","01","01"), 21|22|29 => Pixel_t'("01","01","01"), 19|20|23|24|25|26|28 => Pixel_t'("01","01","10"), 17|18|27 => Pixel_t'("01","10","10"), 1|2|3|4|5|12|13|14|15|16|30|31|32|33|34|35|36|54|55|57 => Pixel_t'("10","10","10"), 6 => Pixel_t'("10","10","11"), 56 => Pixel_t'("10","11","10"), 7|8 => Pixel_t'("10","11","11"), 9|10|11 => Pixel_t'("11","11","11")),
        4 => (0|1|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|32|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","00","01"), 11|31|33|36|52 => Pixel_t'("01","01","01"), 5 => Pixel_t'("01","01","10"), 2|30 => Pixel_t'("01","10","10"), 3|4|6|7|34|35|53|54|55|56|57|58 => Pixel_t'("10","10","10"), 8 => Pixel_t'("10","10","11"), 9|10 => Pixel_t'("11","11","11")),
        5 => (0|1|18|19|20|21|22|23|24|25|26|27|36|37|38|39|40|41|42|43|44|45|46|47|48|49|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 17 => Pixel_t'("00","00","01"), 16|28 => Pixel_t'("00","01","01"), 2|3|11|12|13|14|15|29|30|31|32|50|61 => Pixel_t'("01","01","01"), 51|60 => Pixel_t'("01","10","10"), 4|5|6|7|8|9|10|33|34|35|52|53|54|55|56|57|58|59 => Pixel_t'("10","10","10")),
        6 => (0|1|2|5|6|7|8|9|10|36|37|44|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 3|4|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|39|40|41|43|45|46|47|65|66|67 => Pixel_t'("01","01","01"), 38|42|48|51|52|53|54|55|56|57|58|64 => Pixel_t'("01","10","10"), 49|50|59|60|61|62|63 => Pixel_t'("10","10","10")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|19|28|29|30|31|32|33|34|35|36|37|73 => Pixel_t'("00","00","00"), 26|43|44 => Pixel_t'("00","01","01"), 18|20|21|22|23|24|25|27|38|41|42|45|46|47|48|49|50|51|52|53|54|55|56|57 => Pixel_t'("01","01","01"), 58|72 => Pixel_t'("01","01","10"), 39|40|59|60|61|62|63|64|65|66|67|68|69|70|71 => Pixel_t'("10","10","10")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|26|27|28|29|30|31|32|33|34|35|36|37|38|49|50|51|52|64|67|68|73 => Pixel_t'("00","00","00"), 21|65|70 => Pixel_t'("00","00","01"), 53|66|69 => Pixel_t'("00","01","01"), 22|23|24|25|42|43|44|45|46|47|48|54|55|56|57|58|59|60|61|62|63|71|72 => Pixel_t'("01","01","01"), 39 => Pixel_t'("01","10","01"), 40|41 => Pixel_t'("10","10","10")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|27|28|29|30|31|32|33|34|35|36|37|48|49|50|51|52|53|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 58 => Pixel_t'("00","01","01"), 24|25|26|47|54|57 => Pixel_t'("01","01","01"), 38|39|42|44|45|46|55|56 => Pixel_t'("10","10","10"), 43 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|28|29|30|31|32|33|34|35|36|47|48|49|50|51|52|53|54|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 25|26|27|46|57|58 => Pixel_t'("01","01","01"), 37|42|45|55|56 => Pixel_t'("10","10","10"), 38|44 => Pixel_t'("10","10","11"), 39|43 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
        11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|29|30|31|32|33|34|35|45|46|47|48|49|50|51|52|53|54|55|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 26 => Pixel_t'("00","01","01"), 27|28|56 => Pixel_t'("01","01","01"), 36|38|39|42|43|44 => Pixel_t'("10","10","10"), 37 => Pixel_t'("10","11","11"), 40|41 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|31|32|33|34|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 30|35 => Pixel_t'("00","01","01"), 28|29 => Pixel_t'("01","01","01"), 36|37|38|39|40|42|43 => Pixel_t'("10","10","10"), 41 => Pixel_t'("10","11","11")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|32|33|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29|30|31|34 => Pixel_t'("01","01","01"), 35|36 => Pixel_t'("01","10","10"), 37|38|39|40|41|42|43 => Pixel_t'("10","10","10")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 30|31|32|33|34|35|36|37|38|39|40 => Pixel_t'("01","01","01"), 41|42 => Pixel_t'("01","10","10"), 43 => Pixel_t'("10","10","10")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|30|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","01","01"), 21|22|23|24|31|32|44 => Pixel_t'("01","01","01"), 25|28|43 => Pixel_t'("01","10","10"), 26|27|33|34|35|36|37|38|39|40|41|42 => Pixel_t'("10","10","10")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 20|45 => Pixel_t'("01","01","01"), 43|44 => Pixel_t'("01","10","10"), 29|42 => Pixel_t'("10","10","10"), 21 => Pixel_t'("10","11","10"), 22|23|24|25|26|27|28|30|31|35|36|41 => Pixel_t'("10","11","11"), 32|33|34|37|38|39|40 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 45 => Pixel_t'("01","10","10"), 20|34|35|44 => Pixel_t'("10","10","10"), 22|23|24|25|26|27|28|29|30|31|32|33|36|37|38|43 => Pixel_t'("10","11","11"), 21|39|40|41|42 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 45 => Pixel_t'("01","01","01"), 20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|44 => Pixel_t'("10","10","10"), 40 => Pixel_t'("11","10","10"), 41|42|43 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 23|24|44|45 => Pixel_t'("01","01","01"), 27 => Pixel_t'("01","10","01"), 25|26|28|29|30|31|43 => Pixel_t'("01","10","10"), 32|33|34|35|36|37|38|39|40|42 => Pixel_t'("10","10","10"), 41 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 44 => Pixel_t'("00","01","01"), 27|28|29|30|31|32|33|34|35|36|41|42|43 => Pixel_t'("01","01","01"), 38 => Pixel_t'("01","01","10"), 37|39 => Pixel_t'("01","10","10"), 40 => Pixel_t'("10","10","10")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 34|35|36|37|38|40|41|42|43|44 => Pixel_t'("01","01","01"), 39 => Pixel_t'("01","01","10")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00"), 42 => Pixel_t'("00","00","01"), 41 => Pixel_t'("00","01","01"), 38|39|40|43 => Pixel_t'("01","01","01")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39|40|41|42|43|44|45|46|47|48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|64|65|66|67|68|69|70|71|72|73 => Pixel_t'("00","00","00")));


    -- SCORE --------------------------------------------------------------------------------------------------------------------------

    constant score_9 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|10|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|10|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|13|14 => Pixel_t'("00","00","00"), 9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_8 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_7 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|3|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_6 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 2|3|4|5 => Pixel_t'("11","11","11")),
        2 => (0|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3|4 => Pixel_t'("11","11","11")),
        3 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        11 => (0|4|13|14 => Pixel_t'("00","00","00"), 1|2|3|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|4|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_5 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|11|14 => Pixel_t'("00","00","00"), 1|2|3|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|11|12|14 => Pixel_t'("00","00","00"), 1|2|3|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_4 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 2|3|11|12 => Pixel_t'("11","11","11")),
        2 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|13|14 => Pixel_t'("00","00","00"), 11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_3 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|1|2|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_2 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        15 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00"), 1|2|3 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|11|12|14 => Pixel_t'("00","00","00"), 1|2|3|13 => Pixel_t'("11","11","11")),
        20 => (0|4|5|6|7|8|9|10|11|14 => Pixel_t'("00","00","00"), 1|2|3|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_1 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|2|3|4|5|11|12|13|14 => Pixel_t'("00","00","00"), 6|7|8|9|10 => Pixel_t'("11","11","11")),
        2 => (0|1|2|11|12|13|14 => Pixel_t'("00","00","00"), 3|4|5|6|7|8|9|10 => Pixel_t'("11","11","11")),
        3 => (0|1|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 2|3|4|8|9|10 => Pixel_t'("11","11","11")),
        4 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        5 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        6 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        7 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        8 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        9 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        10 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        11 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        12 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        13 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        14 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        15 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        16 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        17 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        18 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        19 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        20 => (0|1|2|3|4|5|6|7|11|12|13|14 => Pixel_t'("00","00","00"), 8|9|10 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));

    constant score_0 : bit_map_t (0 to score_sizeY-1, 0 to score_sizeX-1) := 
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")),
        1 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        2 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        3 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        4 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        5 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        6 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        7 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        8 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        9 => (0|4|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|10|11|12|13 => Pixel_t'("11","11","11")),
        10 => (0|4|5|6|7|8|10|14 => Pixel_t'("00","00","00"), 1|2|3|9|11|12|13 => Pixel_t'("11","11","11")),
        11 => (0|4|5|6|7|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|8|11|12|13 => Pixel_t'("11","11","11")),
        12 => (0|4|5|6|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|7|11|12|13 => Pixel_t'("11","11","11")),
        13 => (0|4|5|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|6|11|12|13 => Pixel_t'("11","11","11")),
        14 => (0|4|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|5|11|12|13 => Pixel_t'("11","11","11")),
        15 => (0|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|4|11|12|13 => Pixel_t'("11","11","11")),
        16 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        17 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        18 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        19 => (0|4|5|6|7|8|9|10|14 => Pixel_t'("00","00","00"), 1|2|3|11|12|13 => Pixel_t'("11","11","11")),
        20 => (0|5|6|7|8|9|14 => Pixel_t'("00","00","00"), 1|2|3|4|10|11|12|13 => Pixel_t'("11","11","11")),
        21 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        22 => (0|14 => Pixel_t'("00","00","00"), 1|2|3|4|5|6|7|8|9|10|11|12|13 => Pixel_t'("11","11","11")),
        23 => (0|1|13|14 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|9|10|11|12 => Pixel_t'("11","11","11")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14 => Pixel_t'("00","00","00")));





    constant ALIEN_1 : bit_map_t (0 to alien1_sizeY-1, 0 to alien1_sizeX-1) :=
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")),
        1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14|15|16|21|22|23|24 => Pixel_t'("00","01","00"), 17|18|19|20 => Pixel_t'("01","01","01")),
        2 => (0|1|2|3|4|5|6|7|8|9|10|11|12|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 13|23 => Pixel_t'("00","01","00"), 15|16 => Pixel_t'("00","01","01"), 14 => Pixel_t'("01","01","01"), 21|22 => Pixel_t'("01","10","01"), 17|20 => Pixel_t'("01","10","10"), 18|19 => Pixel_t'("10","11","10")),
        3 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17 => Pixel_t'("01","01","01"), 22|24 => Pixel_t'("01","10","01"), 21 => Pixel_t'("01","10","10"), 19|20|23 => Pixel_t'("01","11","10"), 18 => Pixel_t'("10","11","10")),
        4 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 23|25 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 18|19|24 => Pixel_t'("10","11","10")),
        5 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","10","01"), 26 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 19|23|24|25 => Pixel_t'("10","11","10")),
        6 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 28 => Pixel_t'("00","01","00"), 25 => Pixel_t'("01","10","01"), 26|27 => Pixel_t'("01","10","10"), 20|21|22 => Pixel_t'("01","11","10"), 19|23|24 => Pixel_t'("10","11","10")),
        7 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 29 => Pixel_t'("00","01","00"), 26 => Pixel_t'("01","10","01"), 27 => Pixel_t'("01","10","10"), 21|24|25|28 => Pixel_t'("01","11","10"), 19 => Pixel_t'("10","10","10"), 20|22|23 => Pixel_t'("10","11","10")),
        8 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 30 => Pixel_t'("00","01","00"), 19|25|26|27|28|29 => Pixel_t'("01","10","01"), 21|22|23|24 => Pixel_t'("01","11","10"), 20 => Pixel_t'("10","11","10")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 31 => Pixel_t'("00","01","00"), 19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'("01","10","01")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 22|26|32 => Pixel_t'("00","01","00"), 21 => Pixel_t'("00","01","01"), 19|23|24|25|27|28|29 => Pixel_t'("00","10","01"), 17|18|20|30|31 => Pixel_t'("01","10","01")),
        11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 16|19|20|21|23|26|27 => Pixel_t'("00","01","00"), 22|24|25 => Pixel_t'("00","10","00"), 28|29|30|31 => Pixel_t'("00","10","01"), 17|18|32 => Pixel_t'("01","10","01")),
        12 => (0|1|2|3|4|5|6|8|9|10|11|12|13|14|15|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 7|16|18|19|20|21|23|24|25|27|28|29|32|33 => Pixel_t'("00","01","00"), 31 => Pixel_t'("00","01","01"), 22 => Pixel_t'("00","10","00"), 26|30 => Pixel_t'("00","10","01"), 17 => Pixel_t'("01","10","01")),
        13 => (0|1|2|11|12|13|14|15|36|37|38|39 => Pixel_t'("00","00","00"), 3|4|9|10|16|28|29|32 => Pixel_t'("00","01","00"), 35 => Pixel_t'("00","01","01"), 27 => Pixel_t'("00","10","00"), 5|6|7|8|18|19|20|25|26|30|31|33 => Pixel_t'("00","10","01"), 17|21|22|23|24|34 => Pixel_t'("01","10","01")),
        14 => (0|1|9|10|39 => Pixel_t'("00","00","00"), 2|3|4|5|6|7|8|11|13|29|30|31|32|33|34|35|36|37|38 => Pixel_t'("00","01","00"), 12 => Pixel_t'("00","01","01"), 14|15|26|27|28 => Pixel_t'("00","10","01"), 16|17|22|25 => Pixel_t'("01","10","01"), 21 => Pixel_t'("01","10","10"), 18|19|23|24 => Pixel_t'("01","11","10"), 20 => Pixel_t'("10","10","10")),
        15 => (0|1|3|10|11|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 2|4|5|6|7|8|9|12|13|14|15|23|24|25|26|27|28|29|30|31|35 => Pixel_t'("00","01","00"), 16|21 => Pixel_t'("00","10","01"), 17|18|19|20|22 => Pixel_t'("01","10","01")),
        16 => (0|1|2|3|9|10|11|12|13|14|15|16|32|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|5|6|7|8|21|22|23|24|25|26|27|28|29|30|31|33|34 => Pixel_t'("00","01","00"), 20 => Pixel_t'("00","10","00"), 19 => Pixel_t'("00","10","01"), 17|18 => Pixel_t'("01","10","01")),
        17 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 20|21|22|23|24|25|26|27|28|29|30|31|32|33 => Pixel_t'("00","01","00"), 17|18|19 => Pixel_t'("00","10","01")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 16|20|21|22|23|24|25|26|27|28|29|30|31|32 => Pixel_t'("00","01","00"), 19 => Pixel_t'("00","10","00"), 18 => Pixel_t'("01","10","01"), 17 => Pixel_t'("01","11","01")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28|29|30|31 => Pixel_t'("00","01","00"), 17|18 => Pixel_t'("01","10","01")),
        20 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18|19|20|21|22|23|24|25|26|27|28|29|30 => Pixel_t'("00","01","00")),
        21 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","01","00")),
        22 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27|28 => Pixel_t'("00","01","00")),
        23 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25|26|27 => Pixel_t'("00","01","00")),
        24 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25 => Pixel_t'("00","01","00"), 26 => Pixel_t'("00","10","01")),
        25 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19|20|21|22|23|24|25 => Pixel_t'("00","01","00")),
        26 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 18|19|21|22|23|24 => Pixel_t'("00","01","00"), 20 => Pixel_t'("00","10","01")),
        27 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17|18|19|22|23 => Pixel_t'("00","01","00"), 14|21 => Pixel_t'("00","01","01"), 20 => Pixel_t'("00","10","01"), 15|16 => Pixel_t'("01","01","01")),
        28 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|22|23|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17|24 => Pixel_t'("00","01","00"), 14|15|16|18|21 => Pixel_t'("00","01","01"), 19|20 => Pixel_t'("01","01","01")),
        29 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")));

    constant ALIEN_2 : bit_map_t (0 to alien2_sizeY-1, 0 to alien2_sizeX-1) :=
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00")),
        1 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|26|27|28|29 => Pixel_t'("00","00","00"), 16|23|24 => Pixel_t'("00","01","00"), 19 => Pixel_t'("00","01","01"), 18|20|21|22|25 => Pixel_t'("01","01","01"), 17 => Pixel_t'("01","10","10")),
        2 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("00","01","00"), 14 => Pixel_t'("01","01","00"), 16|17|18|19|20|21|22|23|24 => Pixel_t'("01","01","01"), 25 => Pixel_t'("10","10","10")),
        3 => (0|1|2|3|4|5|6|7|8|9|10|11|12|27|28|29 => Pixel_t'("00","00","00"), 13|15|16|17 => Pixel_t'("00","01","00"), 24 => Pixel_t'("00","01","01"), 18|19|20|21|22|23|26 => Pixel_t'("01","01","01"), 14 => Pixel_t'("01","10","01"), 25 => Pixel_t'("10","10","10")),
        4 => (0|1|2|7|8|9|10|11|12|18|19|20|21|22|29 => Pixel_t'("00","00","00"), 3|4|6|16|17|23|24 => Pixel_t'("00","01","00"), 5|13|26|27|28 => Pixel_t'("01","01","01"), 14|15 => Pixel_t'("01","10","01"), 25 => Pixel_t'("01","10","10")),
        5 => (0|1|18|19|20|21|22 => Pixel_t'("00","00","00"), 9|12|13|14|15|16|17|23|24|26|27 => Pixel_t'("00","01","00"), 2|3 => Pixel_t'("01","01","00"), 4|8|10|11|29 => Pixel_t'("01","01","01"), 5|6|7|25|28 => Pixel_t'("01","10","01")),
        6 => (0|14|15|19|20|21|22 => Pixel_t'("00","00","00"), 1|2|3|12|13|16|17|18|29 => Pixel_t'("00","01","00"), 4|5 => Pixel_t'("01","01","00"), 6|7|8|9|11|23|24|25|26|27|28 => Pixel_t'("01","01","01"), 10 => Pixel_t'("01","10","01")),
        7 => (0|1|29 => Pixel_t'("00","00","00"), 2|3|4|5|7|8|9|10|11|12|13|14|15|16|17|28 => Pixel_t'("00","01","00"), 18|19 => Pixel_t'("01","01","01"), 6|20|22|25|26|27 => Pixel_t'("01","10","01"), 21|24 => Pixel_t'("01","10","10"), 23 => Pixel_t'("10","10","10")),
        8 => (0|1|2|3|4|5|7|8|9|10|11|12|13|14|15|16|28|29 => Pixel_t'("00","00","00"), 6|17 => Pixel_t'("00","01","00"), 27 => Pixel_t'("01","01","01"), 18|19|26 => Pixel_t'("01","10","01"), 20|21|23 => Pixel_t'("01","10","10"), 22|24|25 => Pixel_t'("10","10","10")),
        9 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|27|28|29 => Pixel_t'("00","00","00"), 26 => Pixel_t'("01","01","01"), 17|18 => Pixel_t'("01","10","01"), 19|20|21|25 => Pixel_t'("01","10","10"), 22|23|24 => Pixel_t'("10","10","10")),
        10 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|25|26|27|28|29 => Pixel_t'("00","00","00"), 16|24 => Pixel_t'("01","01","01"), 17 => Pixel_t'("01","10","01"), 18|19|20|21|23 => Pixel_t'("01","10","10"), 22 => Pixel_t'("10","10","10")),
        11 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 22 => Pixel_t'("01","01","01"), 16|17 => Pixel_t'("01","10","01"), 18 => Pixel_t'("01","10","10"), 19|20|21 => Pixel_t'("10","10","10")),
        12 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("00","01","00"), 16|17 => Pixel_t'("01","01","01"), 18|20 => Pixel_t'("01","10","01"), 19 => Pixel_t'("10","10","10")),
        13 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15|17|18 => Pixel_t'("01","01","01"), 16 => Pixel_t'("01","10","01")),
        14 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","01","01"), 15|16|17 => Pixel_t'("01","10","01")),
        15 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14 => Pixel_t'("00","01","00"), 18 => Pixel_t'("01","01","01"), 15|16|17 => Pixel_t'("01","10","01")),
        16 => (0|1|2|3|4|5|6|7|8|9|10|11|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 12 => Pixel_t'("00","01","00"), 13|17 => Pixel_t'("01","01","01"), 14|15|16 => Pixel_t'("01","10","01")),
        17 => (0|1|2|3|4|5|6|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14|15|17 => Pixel_t'("00","01","00"), 7|12|13|16 => Pixel_t'("01","01","01"), 8|9|10|11 => Pixel_t'("10","10","10")),
        18 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 14|17 => Pixel_t'("00","01","00"), 15 => Pixel_t'("01","10","01"), 16 => Pixel_t'("10","10","10")),
        19 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|17|18|19|20|21|22|23|24|25|26|27|28|29 => Pixel_t'("00","00","00"), 15 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","10","10")));

    constant ALIEN_3 : bit_map_t (0 to alien3_sizeY-1, 0 to alien3_sizeX-1) :=
        (0 => (0|1|2|7|8|9 => Pixel_t'("00","00","00"), 6 => Pixel_t'("01","01","00"), 3 => Pixel_t'("10","01","00"), 4|5 => Pixel_t'("11","10","00")),
        1 => (0|1|8|9 => Pixel_t'("00","00","00"), 2|7 => Pixel_t'("00","01","00"), 6 => Pixel_t'("01","10","00"), 3|4|5 => Pixel_t'("11","10","00")),
        2 => (0|8|9 => Pixel_t'("00","00","00"), 1|7 => Pixel_t'("00","01","00"), 2 => Pixel_t'("00","10","00"), 3 => Pixel_t'("01","01","00"), 6 => Pixel_t'("01","10","00"), 4|5 => Pixel_t'("10","10","00")),
        3 => (0|3|9 => Pixel_t'("00","00","00"), 4|6|7|8 => Pixel_t'("00","01","00"), 1|2|5 => Pixel_t'("00","10","00")),
        4 => (0|3|9 => Pixel_t'("00","00","00"), 4|6|7|8 => Pixel_t'("00","01","00"), 1|2|5 => Pixel_t'("00","10","00")),
        5 => (0|1|8|9 => Pixel_t'("00","00","00"), 7 => Pixel_t'("00","01","00"), 2 => Pixel_t'("00","10","00"), 4|6 => Pixel_t'("01","10","00"), 3|5 => Pixel_t'("10","10","00")),
        6 => (0|1|8|9 => Pixel_t'("00","00","00"), 3|5|6|7 => Pixel_t'("00","01","00"), 2|4 => Pixel_t'("00","10","00")),
        7 => (0|3|6|9 => Pixel_t'("00","00","00"), 1|2|4|5|7|8 => Pixel_t'("00","01","00")),
        8 => (2|3|6|7 => Pixel_t'("00","00","00"), 0|1|4|5|8|9 => Pixel_t'("00","01","00")),
        9 => (1|2|3|5|6|7|8 => Pixel_t'("00","00","00"), 0|4|9 => Pixel_t'("00","01","00")));

    constant ASTEROID : bit_map_t (0 to asteroid_sizeY-1, 0 to asteroid_sizeX-1) :=
        (0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|15|16|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14|19 => Pixel_t'("00","01","01"), 17|20|21|22|23 => Pixel_t'("01","01","01"), 18 => Pixel_t'("01","01","10")),
        1 => (0|1|2|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 5|9 => Pixel_t'("00","01","01"), 3|4|6|7|8|10|15|16|17|18|19|20|21|23|24|25|28|29|30 => Pixel_t'("01","01","01"), 11 => Pixel_t'("01","10","10"), 33 => Pixel_t'("10","01","01"), 12|13|14|22|26|27|31|32 => Pixel_t'("10","10","10")),
        2 => (0|9|10|11|39 => Pixel_t'("00","00","00"), 4|5|12|15|17|18|19|20|21|22|23|32|33|34|38 => Pixel_t'("01","01","01"), 35 => Pixel_t'("01","01","10"), 13|30 => Pixel_t'("10","01","01"), 1|2|8|14|16|24|27|28|29|31|36|37 => Pixel_t'("10","10","10"), 3|6|7|25|26 => Pixel_t'("11","11","11")),
        3 => (0|5|15|16|28|31|39 => Pixel_t'("00","00","00"), 27 => Pixel_t'("01","00","00"), 1|11|12|14|17|19|20|21|25|26|29|30|32|33|34|35|36|37|38 => Pixel_t'("01","01","01"), 18 => Pixel_t'("10","01","01"), 2|3|4|6|8|9|10|22|23|24 => Pixel_t'("10","10","10"), 7|13 => Pixel_t'("11","11","11")),
        4 => (0|5|25|26|28|30|31|32|36|39 => Pixel_t'("00","00","00"), 34 => Pixel_t'("01","00","00"), 27 => Pixel_t'("01","00","01"), 1|6|16|17|20|21|22|23|24|29|33|35|37|38 => Pixel_t'("01","01","01"), 3|4|11|12|15|18|19 => Pixel_t'("10","10","10"), 2|7|8|9|10|13|14 => Pixel_t'("11","11","11")),
        5 => (0|17|20|21|22|23|24|25|26|27|28|30|31|32|39 => Pixel_t'("00","00","00"), 29|35|36 => Pixel_t'("01","00","00"), 34 => Pixel_t'("01","01","00"), 6|33|37|38 => Pixel_t'("01","01","01"), 1|3|5|7|8|10|16|18 => Pixel_t'("10","10","10"), 2|4|19 => Pixel_t'("11","10","10"), 9|11|12|13|14|15 => Pixel_t'("11","11","11")),
        6 => (0|6|17|21|22|23|24|25|26|27|28|29|34|35|39 => Pixel_t'("00","00","00"), 30|32 => Pixel_t'("01","00","00"), 5|20|31|33|36|37|38 => Pixel_t'("01","01","01"), 1|2|3|4|7|8|9|10|11|13|14|16|18 => Pixel_t'("10","10","10"), 12 => Pixel_t'("11","10","10"), 15|19 => Pixel_t'("11","11","11")),
        7 => (0|17|21|22|23|24|25|26|27|28|29|32|33|34|35|39 => Pixel_t'("00","00","00"), 30|31 => Pixel_t'("01","00","00"), 3|6|11|20|36|37|38 => Pixel_t'("01","01","01"), 1|2|5|7|8|9|10|16|18 => Pixel_t'("10","10","10"), 4|14 => Pixel_t'("11","10","10"), 12|13|15|19 => Pixel_t'("11","11","11")),
        8 => (0|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|39 => Pixel_t'("00","00","00"), 38 => Pixel_t'("00","00","01"), 1|3|5|9|17|20|36|37 => Pixel_t'("01","01","01"), 2|4|6|7|8|10|11|13|14|15|16 => Pixel_t'("10","10","10"), 12|18|19 => Pixel_t'("11","11","11")),
        9 => (0|21|22|23|24|25|26|27|28|29|30|32|33|34|38|39 => Pixel_t'("00","00","00"), 31|35|36 => Pixel_t'("01","00","00"), 1|7|13|14|17|20|37 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","01","01"), 2|3|4|5|6|8|9|10|11 => Pixel_t'("10","10","10"), 12|15|18|19 => Pixel_t'("11","11","11")),
        10 => (0|1|14|21|22|23|24|25|26|27|28|29|32|33|34|38|39 => Pixel_t'("00","00","00"), 30|31 => Pixel_t'("01","00","00"), 6 => Pixel_t'("01","01","00"), 5|7|8|11|13|20|35|36|37 => Pixel_t'("01","01","01"), 10|16 => Pixel_t'("10","01","01"), 2|4|9|17 => Pixel_t'("10","10","10"), 3 => Pixel_t'("11","10","10"), 19 => Pixel_t'("11","11","10"), 12|15|18 => Pixel_t'("11","11","11")),
        11 => (0|1|6|14|21|22|23|24|25|26|27|28|29|30|32|33|38|39 => Pixel_t'("00","00","00"), 5|7|8|11|13|16|20|31|34|35|36|37 => Pixel_t'("01","01","01"), 3 => Pixel_t'("10","10","01"), 2|4|9|10|17 => Pixel_t'("10","10","10"), 15|19 => Pixel_t'("11","10","10"), 12|18 => Pixel_t'("11","11","11")),
        12 => (0|1|3|6|14|21|22|23|24|25|26|27|28|30|31|32|33|38|39 => Pixel_t'("00","00","00"), 29|35 => Pixel_t'("01","00","00"), 2|7|8|13|16|20|34|36|37 => Pixel_t'("01","01","01"), 4|5|9|10|11|15|17|19 => Pixel_t'("10","10","10"), 12|18 => Pixel_t'("11","10","10")),
        13 => (0|3|21|22|23|24|25|26|27|28|29|30|31|32|33|38|39 => Pixel_t'("00","00","00"), 20|35 => Pixel_t'("01","00","00"), 8 => Pixel_t'("01","01","00"), 1|5|6|7|10|14|17|34|36|37 => Pixel_t'("01","01","01"), 4|11|15|16 => Pixel_t'("10","01","01"), 9|12|18|19 => Pixel_t'("10","10","10"), 2|13 => Pixel_t'("11","10","10")),
        14 => (0|3|21|22|23|24|25|26|27|28|29|30|31|32|38|39 => Pixel_t'("00","00","00"), 20|34|35 => Pixel_t'("01","00","00"), 1|4|5|8|11|12|14|17|33|36|37 => Pixel_t'("01","01","01"), 18 => Pixel_t'("10","01","01"), 6|7|9|10|15|16|19 => Pixel_t'("10","10","10"), 13 => Pixel_t'("11","10","10"), 2 => Pixel_t'("11","11","10")),
        15 => (0|1|21|22|23|24|25|26|27|28|29|30|31|32|34|35|37|38|39 => Pixel_t'("00","00","00"), 3 => Pixel_t'("01","01","00"), 4|5|12|14|15|18|20|33|36 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","01","01"), 13|17 => Pixel_t'("10","10","01"), 6|7|8|9|10|11|19 => Pixel_t'("10","10","10"), 2 => Pixel_t'("11","10","10")),
        16 => (0|1|21|22|23|24|25|26|29|30|32|37|38|39 => Pixel_t'("00","00","00"), 27|28|34 => Pixel_t'("01","00","00"), 2|3|5|11|13|19|20|31|33|35|36 => Pixel_t'("01","01","01"), 6|10|15|17 => Pixel_t'("10","01","01"), 14 => Pixel_t'("10","10","01"), 4|7|8|9|12|16|18 => Pixel_t'("10","10","10")),
        17 => (0|1|17|21|22|23|24|25|26|27|29|30|32|38|39 => Pixel_t'("00","00","00"), 37 => Pixel_t'("00","00","01"), 28|31 => Pixel_t'("01","00","00"), 2|3|5|19|20|33|34|35|36 => Pixel_t'("01","01","01"), 6|15 => Pixel_t'("10","01","01"), 8|16|18 => Pixel_t'("10","10","01"), 4|7|9|10|11|12|13|14 => Pixel_t'("10","10","10")),
        18 => (0|1|21|22|23|24|25|26|27|28|29|30|31|35|37|38|39 => Pixel_t'("00","00","00"), 33 => Pixel_t'("00","01","00"), 34 => Pixel_t'("01","00","00"), 20|32 => Pixel_t'("01","01","00"), 2|3|6|7|15|17|18|36 => Pixel_t'("01","01","01"), 14|19 => Pixel_t'("10","01","01"), 8|13 => Pixel_t'("10","10","01"), 4|5|9|10|11|12|16 => Pixel_t'("10","10","10")),
        19 => (0|1|21|22|23|24|25|26|27|28|29|30|34|35|37|38|39 => Pixel_t'("00","00","00"), 33 => Pixel_t'("00","01","00"), 18|20|31 => Pixel_t'("01","00","00"), 32 => Pixel_t'("01","01","00"), 2|3|6|7|10|13|15|19|36 => Pixel_t'("01","01","01"), 11|16 => Pixel_t'("10","01","01"), 4|9|12|17 => Pixel_t'("10","10","01"), 5|8|14 => Pixel_t'("10","10","10")),
        20 => (0|1|10|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","00","00"), 7 => Pixel_t'("01","01","00"), 2|3|6|9|11|12|13|15|16|19|20|36 => Pixel_t'("01","01","01"), 4|5|17 => Pixel_t'("10","01","01"), 8|14 => Pixel_t'("10","10","01")),
        21 => (0|1|7|10|21|22|23|24|25|26|27|28|29|30|31|32|33|34|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","00","00"), 2|4|6|8|9|11|12|13|16|19|20|35|36 => Pixel_t'("01","01","01"), 3|5|14|15|17 => Pixel_t'("10","01","01")),
        22 => (0|1|4|10|21|22|23|24|25|26|27|28|29|30|31|32|33|35|36|37|38|39 => Pixel_t'("00","00","00"), 34 => Pixel_t'("01","00","00"), 6 => Pixel_t'("01","01","00"), 2|5|7|8|9|11|12|13|14|16|18|19|20 => Pixel_t'("01","01","01"), 17 => Pixel_t'("10","01","01"), 15 => Pixel_t'("10","10","01"), 3 => Pixel_t'("10","10","10")),
        23 => (0|1|2|6|10|20|21|22|23|24|25|26|27|28|29|31|32|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|8|13|30 => Pixel_t'("01","00","00"), 7|33 => Pixel_t'("01","01","00"), 5|9|11|14|15|17|18|19 => Pixel_t'("01","01","01"), 12|16 => Pixel_t'("10","01","01"), 3 => Pixel_t'("10","10","10")),
        24 => (0|1|2|7|8|20|21|22|23|24|25|26|27|28|29|31|32|34|35|37|38|39 => Pixel_t'("00","00","00"), 13|17|36 => Pixel_t'("01","00","00"), 33 => Pixel_t'("01","01","00"), 4|6|14|15|16|18|30 => Pixel_t'("01","01","01"), 9|10|19 => Pixel_t'("10","01","01"), 5|11 => Pixel_t'("10","10","01"), 3|12 => Pixel_t'("10","10","10")),
        25 => (0|1|2|8|14|15|17|21|22|23|24|25|26|27|28|29|31|32|33|34|35|37|38|39 => Pixel_t'("00","00","00"), 18|20 => Pixel_t'("01","00","00"), 13|36 => Pixel_t'("01","01","00"), 4|5|6|7|9|16|19|30 => Pixel_t'("01","01","01"), 11 => Pixel_t'("10","10","01"), 3|10|12 => Pixel_t'("10","10","10")),
        26 => (0|1|2|15|18|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 8|14|20 => Pixel_t'("01","00","00"), 4|6|7|13|16|17|19 => Pixel_t'("01","01","01"), 9|11 => Pixel_t'("10","01","01"), 3|5|10|12 => Pixel_t'("10","10","01")),
        27 => (0|1|2|15|21|22|23|24|25|26|27|28|29|30|31|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 18|20 => Pixel_t'("01","00","00"), 8|35 => Pixel_t'("01","01","00"), 4|9|10|13|14|16|17|19 => Pixel_t'("01","01","01"), 3|7|11|12 => Pixel_t'("10","01","01"), 5|6 => Pixel_t'("10","10","10")),
        28 => (0|1|2|9|15|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 35 => Pixel_t'("01","00","00"), 3|6|10|13|16|17|18|19 => Pixel_t'("01","01","01"), 4|7|11|12|14 => Pixel_t'("10","01","01"), 5 => Pixel_t'("10","10","01"), 8 => Pixel_t'("10","10","10")),
        29 => (0|1|2|3|15|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|7 => Pixel_t'("01","00","00"), 9|13|18 => Pixel_t'("01","01","00"), 6|10|12|14|16|17|19 => Pixel_t'("01","01","01"), 5|8|11 => Pixel_t'("10","01","01")),
        30 => (0|1|2|3|4|5|7|13|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 12|16 => Pixel_t'("01","01","00"), 6|8|10|11|14|17|19 => Pixel_t'("01","01","01"), 9 => Pixel_t'("10","10","01")),
        31 => (0|1|2|3|4|5|6|7|14|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 8|15 => Pixel_t'("01","00","00"), 12|13 => Pixel_t'("01","01","00"), 10|11|17|19 => Pixel_t'("01","01","01"), 9|16 => Pixel_t'("10","01","01")),
        32 => (0|1|2|3|4|5|6|7|8|14|15|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 9 => Pixel_t'("01","00","00"), 10|11|13|16|17 => Pixel_t'("01","01","01"), 12 => Pixel_t'("10","01","01")),
        33 => (0|1|2|3|4|5|6|7|8|9|10|15|18|19|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 20 => Pixel_t'("01","00","00"), 13|14|16 => Pixel_t'("01","01","00"), 11|12|17 => Pixel_t'("01","01","01")),
        34 => (0|1|2|3|4|5|6|7|8|9|10|11|12|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 13 => Pixel_t'("01","00","00"), 14 => Pixel_t'("01","01","00"), 16|17|19 => Pixel_t'("01","01","01")),
        35 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14 => Pixel_t'("01","01","00"), 16|17|19 => Pixel_t'("01","01","01")),
        36 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19 => Pixel_t'("01","01","00"), 16|17 => Pixel_t'("01","01","01")),
        37 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17 => Pixel_t'("01","00","00"), 19 => Pixel_t'("01","01","01")),
        38 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19 => Pixel_t'("01","01","00")),
        39 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")));


end package;