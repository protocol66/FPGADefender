(0 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|15|16|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14|19 => Pixel_t'("00","01","01"), 17|20|21|22|23 => Pixel_t'("01","01","01"), 18 => Pixel_t'("01","01","10")),
1 => (0|1|2|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 5|9 => Pixel_t'("00","01","01"), 3|4|6|7|8|10|15|16|17|18|19|20|21|23|24|25|28|29|30 => Pixel_t'("01","01","01"), 11 => Pixel_t'("01","10","10"), 33 => Pixel_t'("10","01","01"), 12|13|14|22|26|27|31|32 => Pixel_t'("10","10","10")),
2 => (0|9|10|11|39 => Pixel_t'("00","00","00"), 4|5|12|15|17|18|19|20|21|22|23|32|33|34|38 => Pixel_t'("01","01","01"), 35 => Pixel_t'("01","01","10"), 13|30 => Pixel_t'("10","01","01"), 1|2|8|14|16|24|27|28|29|31|36|37 => Pixel_t'("10","10","10"), 3|6|7|25|26 => Pixel_t'("11","11","11")),
3 => (0|5|15|16|28|31|39 => Pixel_t'("00","00","00"), 27 => Pixel_t'("01","00","00"), 1|11|12|14|17|19|20|21|25|26|29|30|32|33|34|35|36|37|38 => Pixel_t'("01","01","01"), 18 => Pixel_t'("10","01","01"), 2|3|4|6|8|9|10|22|23|24 => Pixel_t'("10","10","10"), 7|13 => Pixel_t'("11","11","11")),
4 => (0|5|25|26|28|30|31|32|36|39 => Pixel_t'("00","00","00"), 34 => Pixel_t'("01","00","00"), 27 => Pixel_t'("01","00","01"), 1|6|16|17|20|21|22|23|24|29|33|35|37|38 => Pixel_t'("01","01","01"), 3|4|11|12|15|18|19 => Pixel_t'("10","10","10"), 2|7|8|9|10|13|14 => Pixel_t'("11","11","11")),
5 => (0|17|20|21|22|23|24|25|26|27|28|30|31|32|39 => Pixel_t'("00","00","00"), 29|35|36 => Pixel_t'("01","00","00"), 34 => Pixel_t'("01","01","00"), 6|33|37|38 => Pixel_t'("01","01","01"), 1|3|5|7|8|10|16|18 => Pixel_t'("10","10","10"), 2|4|19 => Pixel_t'("11","10","10"), 9|11|12|13|14|15 => Pixel_t'("11","11","11")),
6 => (0|6|17|21|22|23|24|25|26|27|28|29|34|35|39 => Pixel_t'("00","00","00"), 30|32 => Pixel_t'("01","00","00"), 5|20|31|33|36|37|38 => Pixel_t'("01","01","01"), 1|2|3|4|7|8|9|10|11|13|14|16|18 => Pixel_t'("10","10","10"), 12 => Pixel_t'("11","10","10"), 15|19 => Pixel_t'("11","11","11")),
7 => (0|17|21|22|23|24|25|26|27|28|29|32|33|34|35|39 => Pixel_t'("00","00","00"), 30|31 => Pixel_t'("01","00","00"), 3|6|11|20|36|37|38 => Pixel_t'("01","01","01"), 1|2|5|7|8|9|10|16|18 => Pixel_t'("10","10","10"), 4|14 => Pixel_t'("11","10","10"), 12|13|15|19 => Pixel_t'("11","11","11")),
8 => (0|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|39 => Pixel_t'("00","00","00"), 38 => Pixel_t'("00","00","01"), 1|3|5|9|17|20|36|37 => Pixel_t'("01","01","01"), 2|4|6|7|8|10|11|13|14|15|16 => Pixel_t'("10","10","10"), 12|18|19 => Pixel_t'("11","11","11")),
9 => (0|21|22|23|24|25|26|27|28|29|30|32|33|34|38|39 => Pixel_t'("00","00","00"), 31|35|36 => Pixel_t'("01","00","00"), 1|7|13|14|17|20|37 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","01","01"), 2|3|4|5|6|8|9|10|11 => Pixel_t'("10","10","10"), 12|15|18|19 => Pixel_t'("11","11","11")),
10 => (0|1|14|21|22|23|24|25|26|27|28|29|32|33|34|38|39 => Pixel_t'("00","00","00"), 30|31 => Pixel_t'("01","00","00"), 6 => Pixel_t'("01","01","00"), 5|7|8|11|13|20|35|36|37 => Pixel_t'("01","01","01"), 10|16 => Pixel_t'("10","01","01"), 2|4|9|17 => Pixel_t'("10","10","10"), 3 => Pixel_t'("11","10","10"), 19 => Pixel_t'("11","11","10"), 12|15|18 => Pixel_t'("11","11","11")),
11 => (0|1|6|14|21|22|23|24|25|26|27|28|29|30|32|33|38|39 => Pixel_t'("00","00","00"), 5|7|8|11|13|16|20|31|34|35|36|37 => Pixel_t'("01","01","01"), 3 => Pixel_t'("10","10","01"), 2|4|9|10|17 => Pixel_t'("10","10","10"), 15|19 => Pixel_t'("11","10","10"), 12|18 => Pixel_t'("11","11","11")),
12 => (0|1|3|6|14|21|22|23|24|25|26|27|28|30|31|32|33|38|39 => Pixel_t'("00","00","00"), 29|35 => Pixel_t'("01","00","00"), 2|7|8|13|16|20|34|36|37 => Pixel_t'("01","01","01"), 4|5|9|10|11|15|17|19 => Pixel_t'("10","10","10"), 12|18 => Pixel_t'("11","10","10")),
13 => (0|3|21|22|23|24|25|26|27|28|29|30|31|32|33|38|39 => Pixel_t'("00","00","00"), 20|35 => Pixel_t'("01","00","00"), 8 => Pixel_t'("01","01","00"), 1|5|6|7|10|14|17|34|36|37 => Pixel_t'("01","01","01"), 4|11|15|16 => Pixel_t'("10","01","01"), 9|12|18|19 => Pixel_t'("10","10","10"), 2|13 => Pixel_t'("11","10","10")),
14 => (0|3|21|22|23|24|25|26|27|28|29|30|31|32|38|39 => Pixel_t'("00","00","00"), 20|34|35 => Pixel_t'("01","00","00"), 1|4|5|8|11|12|14|17|33|36|37 => Pixel_t'("01","01","01"), 18 => Pixel_t'("10","01","01"), 6|7|9|10|15|16|19 => Pixel_t'("10","10","10"), 13 => Pixel_t'("11","10","10"), 2 => Pixel_t'("11","11","10")),
15 => (0|1|21|22|23|24|25|26|27|28|29|30|31|32|34|35|37|38|39 => Pixel_t'("00","00","00"), 3 => Pixel_t'("01","01","00"), 4|5|12|14|15|18|20|33|36 => Pixel_t'("01","01","01"), 16 => Pixel_t'("10","01","01"), 13|17 => Pixel_t'("10","10","01"), 6|7|8|9|10|11|19 => Pixel_t'("10","10","10"), 2 => Pixel_t'("11","10","10")),
16 => (0|1|21|22|23|24|25|26|29|30|32|37|38|39 => Pixel_t'("00","00","00"), 27|28|34 => Pixel_t'("01","00","00"), 2|3|5|11|13|19|20|31|33|35|36 => Pixel_t'("01","01","01"), 6|10|15|17 => Pixel_t'("10","01","01"), 14 => Pixel_t'("10","10","01"), 4|7|8|9|12|16|18 => Pixel_t'("10","10","10")),
17 => (0|1|17|21|22|23|24|25|26|27|29|30|32|38|39 => Pixel_t'("00","00","00"), 37 => Pixel_t'("00","00","01"), 28|31 => Pixel_t'("01","00","00"), 2|3|5|19|20|33|34|35|36 => Pixel_t'("01","01","01"), 6|15 => Pixel_t'("10","01","01"), 8|16|18 => Pixel_t'("10","10","01"), 4|7|9|10|11|12|13|14 => Pixel_t'("10","10","10")),
18 => (0|1|21|22|23|24|25|26|27|28|29|30|31|35|37|38|39 => Pixel_t'("00","00","00"), 33 => Pixel_t'("00","01","00"), 34 => Pixel_t'("01","00","00"), 20|32 => Pixel_t'("01","01","00"), 2|3|6|7|15|17|18|36 => Pixel_t'("01","01","01"), 14|19 => Pixel_t'("10","01","01"), 8|13 => Pixel_t'("10","10","01"), 4|5|9|10|11|12|16 => Pixel_t'("10","10","10")),
19 => (0|1|21|22|23|24|25|26|27|28|29|30|34|35|37|38|39 => Pixel_t'("00","00","00"), 33 => Pixel_t'("00","01","00"), 18|20|31 => Pixel_t'("01","00","00"), 32 => Pixel_t'("01","01","00"), 2|3|6|7|10|13|15|19|36 => Pixel_t'("01","01","01"), 11|16 => Pixel_t'("10","01","01"), 4|9|12|17 => Pixel_t'("10","10","01"), 5|8|14 => Pixel_t'("10","10","10")),
20 => (0|1|10|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","00","00"), 7 => Pixel_t'("01","01","00"), 2|3|6|9|11|12|13|15|16|19|20|36 => Pixel_t'("01","01","01"), 4|5|17 => Pixel_t'("10","01","01"), 8|14 => Pixel_t'("10","10","01")),
21 => (0|1|7|10|21|22|23|24|25|26|27|28|29|30|31|32|33|34|37|38|39 => Pixel_t'("00","00","00"), 18 => Pixel_t'("01","00","00"), 2|4|6|8|9|11|12|13|16|19|20|35|36 => Pixel_t'("01","01","01"), 3|5|14|15|17 => Pixel_t'("10","01","01")),
22 => (0|1|4|10|21|22|23|24|25|26|27|28|29|30|31|32|33|35|36|37|38|39 => Pixel_t'("00","00","00"), 34 => Pixel_t'("01","00","00"), 6 => Pixel_t'("01","01","00"), 2|5|7|8|9|11|12|13|14|16|18|19|20 => Pixel_t'("01","01","01"), 17 => Pixel_t'("10","01","01"), 15 => Pixel_t'("10","10","01"), 3 => Pixel_t'("10","10","10")),
23 => (0|1|2|6|10|20|21|22|23|24|25|26|27|28|29|31|32|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|8|13|30 => Pixel_t'("01","00","00"), 7|33 => Pixel_t'("01","01","00"), 5|9|11|14|15|17|18|19 => Pixel_t'("01","01","01"), 12|16 => Pixel_t'("10","01","01"), 3 => Pixel_t'("10","10","10")),
24 => (0|1|2|7|8|20|21|22|23|24|25|26|27|28|29|31|32|34|35|37|38|39 => Pixel_t'("00","00","00"), 13|17|36 => Pixel_t'("01","00","00"), 33 => Pixel_t'("01","01","00"), 4|6|14|15|16|18|30 => Pixel_t'("01","01","01"), 9|10|19 => Pixel_t'("10","01","01"), 5|11 => Pixel_t'("10","10","01"), 3|12 => Pixel_t'("10","10","10")),
25 => (0|1|2|8|14|15|17|21|22|23|24|25|26|27|28|29|31|32|33|34|35|37|38|39 => Pixel_t'("00","00","00"), 18|20 => Pixel_t'("01","00","00"), 13|36 => Pixel_t'("01","01","00"), 4|5|6|7|9|16|19|30 => Pixel_t'("01","01","01"), 11 => Pixel_t'("10","10","01"), 3|10|12 => Pixel_t'("10","10","10")),
26 => (0|1|2|15|18|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 8|14|20 => Pixel_t'("01","00","00"), 4|6|7|13|16|17|19 => Pixel_t'("01","01","01"), 9|11 => Pixel_t'("10","01","01"), 3|5|10|12 => Pixel_t'("10","10","01")),
27 => (0|1|2|15|21|22|23|24|25|26|27|28|29|30|31|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 18|20 => Pixel_t'("01","00","00"), 8|35 => Pixel_t'("01","01","00"), 4|9|10|13|14|16|17|19 => Pixel_t'("01","01","01"), 3|7|11|12 => Pixel_t'("10","01","01"), 5|6 => Pixel_t'("10","10","10")),
28 => (0|1|2|9|15|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|36|37|38|39 => Pixel_t'("00","00","00"), 35 => Pixel_t'("01","00","00"), 3|6|10|13|16|17|18|19 => Pixel_t'("01","01","01"), 4|7|11|12|14 => Pixel_t'("10","01","01"), 5 => Pixel_t'("10","10","01"), 8 => Pixel_t'("10","10","10")),
29 => (0|1|2|3|15|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 4|7 => Pixel_t'("01","00","00"), 9|13|18 => Pixel_t'("01","01","00"), 6|10|12|14|16|17|19 => Pixel_t'("01","01","01"), 5|8|11 => Pixel_t'("10","01","01")),
30 => (0|1|2|3|4|5|7|13|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 12|16 => Pixel_t'("01","01","00"), 6|8|10|11|14|17|19 => Pixel_t'("01","01","01"), 9 => Pixel_t'("10","10","01")),
31 => (0|1|2|3|4|5|6|7|14|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 8|15 => Pixel_t'("01","00","00"), 12|13 => Pixel_t'("01","01","00"), 10|11|17|19 => Pixel_t'("01","01","01"), 9|16 => Pixel_t'("10","01","01")),
32 => (0|1|2|3|4|5|6|7|8|14|15|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 9 => Pixel_t'("01","00","00"), 10|11|13|16|17 => Pixel_t'("01","01","01"), 12 => Pixel_t'("10","01","01")),
33 => (0|1|2|3|4|5|6|7|8|9|10|15|18|19|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 20 => Pixel_t'("01","00","00"), 13|14|16 => Pixel_t'("01","01","00"), 11|12|17 => Pixel_t'("01","01","01")),
34 => (0|1|2|3|4|5|6|7|8|9|10|11|12|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 13 => Pixel_t'("01","00","00"), 14 => Pixel_t'("01","01","00"), 16|17|19 => Pixel_t'("01","01","01")),
35 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 14 => Pixel_t'("01","01","00"), 16|17|19 => Pixel_t'("01","01","01")),
36 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19 => Pixel_t'("01","01","00"), 16|17 => Pixel_t'("01","01","01")),
37 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 17 => Pixel_t'("01","00","00"), 19 => Pixel_t'("01","01","01")),
38 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00"), 19 => Pixel_t'("01","01","00")),
39 => (0|1|2|3|4|5|6|7|8|9|10|11|12|13|14|15|16|17|18|19|20|21|22|23|24|25|26|27|28|29|30|31|32|33|34|35|36|37|38|39 => Pixel_t'("00","00","00")));