(0 => (0|1|2|7|8|9 => Pixel_t'("00","00","00"), 6 => Pixel_t'("01","01","00"), 3 => Pixel_t'("10","01","00"), 4|5 => Pixel_t'("11","10","00")),
1 => (0|1|8|9 => Pixel_t'("00","00","00"), 2|7 => Pixel_t'("00","01","00"), 6 => Pixel_t'("01","10","00"), 3|4|5 => Pixel_t'("11","10","00")),
2 => (0|8|9 => Pixel_t'("00","00","00"), 1|7 => Pixel_t'("00","01","00"), 2 => Pixel_t'("00","10","00"), 3 => Pixel_t'("01","01","00"), 6 => Pixel_t'("01","10","00"), 4|5 => Pixel_t'("10","10","00")),
3 => (0|3|9 => Pixel_t'("00","00","00"), 4|6|7|8 => Pixel_t'("00","01","00"), 1|2|5 => Pixel_t'("00","10","00")),
4 => (0|3|9 => Pixel_t'("00","00","00"), 4|6|7|8 => Pixel_t'("00","01","00"), 1|2|5 => Pixel_t'("00","10","00")),
5 => (0|1|8|9 => Pixel_t'("00","00","00"), 7 => Pixel_t'("00","01","00"), 2 => Pixel_t'("00","10","00"), 4|6 => Pixel_t'("01","10","00"), 3|5 => Pixel_t'("10","10","00")),
6 => (0|1|8|9 => Pixel_t'("00","00","00"), 3|5|6|7 => Pixel_t'("00","01","00"), 2|4 => Pixel_t'("00","10","00")),
7 => (0|3|6|9 => Pixel_t'("00","00","00"), 1|2|4|5|7|8 => Pixel_t'("00","01","00")),
8 => (2|3|6|7 => Pixel_t'("00","00","00"), 0|1|4|5|8|9 => Pixel_t'("00","01","00")),
9 => (1|2|3|5|6|7|8 => Pixel_t'("00","00","00"), 0|4|9 => Pixel_t'("00","01","00")));