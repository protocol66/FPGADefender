library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.my_data_types.all;

package bitmaps is
    constant BACKGROUND : Pixel_t := BLACK;

    constant DEFUALT_OBJ : OBJ := (box => Bounding_Box'(0,0,0,0,'0', 1, 1), 
                                   bit_map => bit_map_t'(0, 0, 1, 1), 
                                   abs_mem_addr => (others=>'0'),
                                   enable => '0', 
                                   in_bounds => '0', 
                                   pixel => BACKGROUND);

    -- These are generated by the img2rom.py script in the utils folder
    constant NULL_BITMAP : bit_map_t := bit_map_t'(0, 0, 1, 1);
    constant LINE_BITMAP : bit_map_t := bit_map_t'(0, 1, 640, 2);
    constant SHIP_BITMAP : bit_map_t := bit_map_t'(0, 1281, 74, 25);
    constant LASER_BITMAP : bit_map_t := bit_map_t'(0, 3131, 12, 3);
    constant SCORE_0_BITMAP : bit_map_t := bit_map_t'(0, 3167, 15, 25);
    constant SCORE_1_BITMAP : bit_map_t := bit_map_t'(0, 3542, 15, 25);
    constant SCORE_2_BITMAP : bit_map_t := bit_map_t'(0, 3917, 15, 25);
    constant SCORE_3_BITMAP : bit_map_t := bit_map_t'(0, 4292, 15, 25);
    constant SCORE_4_BITMAP : bit_map_t := bit_map_t'(0, 4667, 15, 25);
    constant SCORE_5_BITMAP : bit_map_t := bit_map_t'(0, 5042, 15, 25);
    constant SCORE_6_BITMAP : bit_map_t := bit_map_t'(0, 5417, 15, 25);
    constant SCORE_7_BITMAP : bit_map_t := bit_map_t'(0, 5792, 15, 25);
    constant SCORE_8_BITMAP : bit_map_t := bit_map_t'(0, 6167, 15, 25);
    constant SCORE_9_BITMAP : bit_map_t := bit_map_t'(0, 6542, 15, 25);
    constant ALIEN1_BITMAP : bit_map_t := bit_map_t'(0, 6917, 39, 30);
    constant ALIEN2_BITMAP : bit_map_t := bit_map_t'(0, 8087, 28, 12);
    constant ALIEN3_BITMAP : bit_map_t := bit_map_t'(0, 8423, 20, 13);
    constant ASTEROID_BITMAP : bit_map_t := bit_map_t'(0, 8683, 40, 40);
    constant START_BITMAP : bit_map_t := bit_map_t'(0, 10283, 250, 100);
    constant GAME_OVER_BITMAP : bit_map_t := bit_map_t'(0, 35283, 380, 73);
    
    
    
                                   

    constant fx1 : Sound_FX_t := (18, (550, 404, 315, 494, 182, 260, 455, 387, 340, 550, 404, 315, 494, 182, 260, 455, 387, 340, others => 0));
    constant fx2 : Sound_FX_t := (10, (300, 350, 500, 700, 990, 970, 1050, 1010, 950, 800, 770, 640, 500, 350, 355, others => 0));
    constant fx3 : Sound_FX_t := (6,  (500, 790, 950, 1300, 1710, 1650, 1300, 800, 700, others=> 0));
    constant fx4 : Sound_FX_t := (60, (1300, 1650, 1660, 1510, 1309, 1158, 1007, 855, others=> 0));
    constant fx5 : Sound_FX_t := (25, (300, 210, 310, 170, 250, 210, 310, 120, 220, 170, 160, 90, 290, 230, 140, 320, 200, 100, 250, 290, others => 0));
    constant fx6 : Sound_FX_t := (15, (700, 702, 698, 701, 699, 700, 250, 251, 249, 252, 248, 130, 131, 129, 132, 128, 130, 130, others=>0));

    -- these constants are legacy support
    constant ship_sizeX : positive := SHIP_BITMAP.x_size;
    constant ship_sizeY : positive := SHIP_BITMAP.y_size;

end package;