../../components/bin2dec.vhdl